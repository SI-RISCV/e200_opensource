 /*                                                                      
 Copyright 2018 Nuclei System Technology, Inc.                
                                                                         
 Licensed under the Apache License, Version 2.0 (the "License");         
 you may not use this file except in compliance with the License.        
 You may obtain a copy of the License at                                 
                                                                         
     http://www.apache.org/licenses/LICENSE-2.0                          
                                                                         
  Unless required by applicable law or agreed to in writing, software    
 distributed under the License is distributed on an "AS IS" BASIS,       
 WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 See the License for the specific language governing permissions and     
 limitations under the License.                                          
 */                                                                      
                                                                         
                                                                         
                                                                         

module sirv_qspi_1cs(
  input   clock,
  input   reset,
  output  io_port_sck,
  input   io_port_dq_0_i,
  output  io_port_dq_0_o,
  output  io_port_dq_0_oe,
  input   io_port_dq_1_i,
  output  io_port_dq_1_o,
  output  io_port_dq_1_oe,
  input   io_port_dq_2_i,
  output  io_port_dq_2_o,
  output  io_port_dq_2_oe,
  input   io_port_dq_3_i,
  output  io_port_dq_3_o,
  output  io_port_dq_3_oe,
  output  io_port_cs_0,
  output  io_tl_i_0_0,
  output  io_tl_r_0_a_ready,
  input   io_tl_r_0_a_valid,
  input  [2:0] io_tl_r_0_a_bits_opcode,
  input  [2:0] io_tl_r_0_a_bits_param,
  input  [2:0] io_tl_r_0_a_bits_size,
  input  [4:0] io_tl_r_0_a_bits_source,
  input  [28:0] io_tl_r_0_a_bits_address,
  input  [3:0] io_tl_r_0_a_bits_mask,
  input  [31:0] io_tl_r_0_a_bits_data,
  input   io_tl_r_0_b_ready,
  output  io_tl_r_0_b_valid,
  output [2:0] io_tl_r_0_b_bits_opcode,
  output [1:0] io_tl_r_0_b_bits_param,
  output [2:0] io_tl_r_0_b_bits_size,
  output [4:0] io_tl_r_0_b_bits_source,
  output [28:0] io_tl_r_0_b_bits_address,
  output [3:0] io_tl_r_0_b_bits_mask,
  output [31:0] io_tl_r_0_b_bits_data,
  output  io_tl_r_0_c_ready,
  input   io_tl_r_0_c_valid,
  input  [2:0] io_tl_r_0_c_bits_opcode,
  input  [2:0] io_tl_r_0_c_bits_param,
  input  [2:0] io_tl_r_0_c_bits_size,
  input  [4:0] io_tl_r_0_c_bits_source,
  input  [28:0] io_tl_r_0_c_bits_address,
  input  [31:0] io_tl_r_0_c_bits_data,
  input   io_tl_r_0_c_bits_error,
  input   io_tl_r_0_d_ready,
  output  io_tl_r_0_d_valid,
  output [2:0] io_tl_r_0_d_bits_opcode,
  output [1:0] io_tl_r_0_d_bits_param,
  output [2:0] io_tl_r_0_d_bits_size,
  output [4:0] io_tl_r_0_d_bits_source,
  output  io_tl_r_0_d_bits_sink,
  output [1:0] io_tl_r_0_d_bits_addr_lo,
  output [31:0] io_tl_r_0_d_bits_data,
  output  io_tl_r_0_d_bits_error,
  output  io_tl_r_0_e_ready,
  input   io_tl_r_0_e_valid,
  input   io_tl_r_0_e_bits_sink
);
  wire [1:0] T_955_fmt_proto;
  wire  T_955_fmt_endian;
  wire  T_955_fmt_iodir;
  wire [3:0] T_955_fmt_len;
  wire [11:0] T_955_sck_div;
  wire  T_955_sck_pol;
  wire  T_955_sck_pha;
  wire  T_955_cs_id;
  wire  T_955_cs_dflt_0;
  wire [1:0] T_955_cs_mode;
  wire [7:0] T_955_dla_cssck;
  wire [7:0] T_955_dla_sckcs;
  wire [7:0] T_955_dla_intercs;
  wire [7:0] T_955_dla_interxfr;
  wire [3:0] T_955_wm_tx;
  wire [3:0] T_955_wm_rx;
  reg [1:0] ctrl_fmt_proto;
  reg [31:0] GEN_236;
  reg  ctrl_fmt_endian;
  reg [31:0] GEN_237;
  reg  ctrl_fmt_iodir;
  reg [31:0] GEN_238;
  reg [3:0] ctrl_fmt_len;
  reg [31:0] GEN_239;
  reg [11:0] ctrl_sck_div;
  reg [31:0] GEN_240;
  reg  ctrl_sck_pol;
  reg [31:0] GEN_241;
  reg  ctrl_sck_pha;
  reg [31:0] GEN_242;
  reg  ctrl_cs_id;
  reg [31:0] GEN_243;
  reg  ctrl_cs_dflt_0;
  reg [31:0] GEN_244;
  reg [1:0] ctrl_cs_mode;
  reg [31:0] GEN_245;
  reg [7:0] ctrl_dla_cssck;
  reg [31:0] GEN_246;
  reg [7:0] ctrl_dla_sckcs;
  reg [31:0] GEN_247;
  reg [7:0] ctrl_dla_intercs;
  reg [31:0] GEN_248;
  reg [7:0] ctrl_dla_interxfr;
  reg [31:0] GEN_249;
  reg [3:0] ctrl_wm_tx;
  reg [31:0] GEN_250;
  reg [3:0] ctrl_wm_rx;
  reg [31:0] GEN_251;
  wire  fifo_clock;
  wire  fifo_reset;
  wire [1:0] fifo_io_ctrl_fmt_proto;
  wire  fifo_io_ctrl_fmt_endian;
  wire  fifo_io_ctrl_fmt_iodir;
  wire [3:0] fifo_io_ctrl_fmt_len;
  wire [1:0] fifo_io_ctrl_cs_mode;
  wire [3:0] fifo_io_ctrl_wm_tx;
  wire [3:0] fifo_io_ctrl_wm_rx;
  wire  fifo_io_link_tx_ready;
  wire  fifo_io_link_tx_valid;
  wire [7:0] fifo_io_link_tx_bits;
  wire  fifo_io_link_rx_valid;
  wire [7:0] fifo_io_link_rx_bits;
  wire [7:0] fifo_io_link_cnt;
  wire [1:0] fifo_io_link_fmt_proto;
  wire  fifo_io_link_fmt_endian;
  wire  fifo_io_link_fmt_iodir;
  wire  fifo_io_link_cs_set;
  wire  fifo_io_link_cs_clear;
  wire  fifo_io_link_cs_hold;
  wire  fifo_io_link_active;
  wire  fifo_io_link_lock;
  wire  fifo_io_tx_ready;
  wire  fifo_io_tx_valid;
  wire [7:0] fifo_io_tx_bits;
  wire  fifo_io_rx_ready;
  wire  fifo_io_rx_valid;
  wire [7:0] fifo_io_rx_bits;
  wire  fifo_io_ip_txwm;
  wire  fifo_io_ip_rxwm;
  wire  mac_clock;
  wire  mac_reset;
  wire  mac_io_port_sck;
  wire  mac_io_port_dq_0_i;
  wire  mac_io_port_dq_0_o;
  wire  mac_io_port_dq_0_oe;
  wire  mac_io_port_dq_1_i;
  wire  mac_io_port_dq_1_o;
  wire  mac_io_port_dq_1_oe;
  wire  mac_io_port_dq_2_i;
  wire  mac_io_port_dq_2_o;
  wire  mac_io_port_dq_2_oe;
  wire  mac_io_port_dq_3_i;
  wire  mac_io_port_dq_3_o;
  wire  mac_io_port_dq_3_oe;
  wire  mac_io_port_cs_0;
  wire [11:0] mac_io_ctrl_sck_div;
  wire  mac_io_ctrl_sck_pol;
  wire  mac_io_ctrl_sck_pha;
  wire [7:0] mac_io_ctrl_dla_cssck;
  wire [7:0] mac_io_ctrl_dla_sckcs;
  wire [7:0] mac_io_ctrl_dla_intercs;
  wire [7:0] mac_io_ctrl_dla_interxfr;
  wire  mac_io_ctrl_cs_id;
  wire  mac_io_ctrl_cs_dflt_0;
  wire  mac_io_link_tx_ready;
  wire  mac_io_link_tx_valid;
  wire [7:0] mac_io_link_tx_bits;
  wire  mac_io_link_rx_valid;
  wire [7:0] mac_io_link_rx_bits;
  wire [7:0] mac_io_link_cnt;
  wire [1:0] mac_io_link_fmt_proto;
  wire  mac_io_link_fmt_endian;
  wire  mac_io_link_fmt_iodir;
  wire  mac_io_link_cs_set;
  wire  mac_io_link_cs_clear;
  wire  mac_io_link_cs_hold;
  wire  mac_io_link_active;
  wire  T_1021_txwm;
  wire  T_1021_rxwm;
  wire [1:0] T_1025;
  wire  T_1026;
  wire  T_1027;
  reg  ie_txwm;
  reg [31:0] GEN_252;
  reg  ie_rxwm;
  reg [31:0] GEN_253;
  wire  T_1030;
  wire  T_1031;
  wire  T_1032;
  wire  T_1036;
  wire  T_1039;
  wire  T_1063_ready;
  wire  T_1063_valid;
  wire  T_1063_bits_read;
  wire [9:0] T_1063_bits_index;
  wire [31:0] T_1063_bits_data;
  wire [3:0] T_1063_bits_mask;
  wire [9:0] T_1063_bits_extra;
  wire  T_1080;
  wire [26:0] T_1081;
  wire [1:0] T_1082;
  wire [6:0] T_1083;
  wire [9:0] T_1084;
  wire  T_1102_ready;
  wire  T_1102_valid;
  wire  T_1102_bits_read;
  wire [31:0] T_1102_bits_data;
  wire [9:0] T_1102_bits_extra;
  wire  T_1138_ready;
  wire  T_1138_valid;
  wire  T_1138_bits_read;
  wire [9:0] T_1138_bits_index;
  wire [31:0] T_1138_bits_data;
  wire [3:0] T_1138_bits_mask;
  wire [9:0] T_1138_bits_extra;
  wire [9:0] T_1223;
  wire  T_1225;
  wire [9:0] T_1231;
  wire [9:0] T_1232;
  wire  T_1234;
  wire [9:0] T_1240;
  wire [9:0] T_1241;
  wire  T_1243;
  wire [9:0] T_1249;
  wire [9:0] T_1250;
  wire  T_1252;
  wire [9:0] T_1258;
  wire [9:0] T_1259;
  wire  T_1261;
  wire [9:0] T_1267;
  wire [9:0] T_1268;
  wire  T_1270;
  wire [9:0] T_1276;
  wire [9:0] T_1277;
  wire  T_1279;
  wire [9:0] T_1285;
  wire [9:0] T_1286;
  wire  T_1288;
  wire [9:0] T_1294;
  wire [9:0] T_1295;
  wire  T_1297;
  wire [9:0] T_1303;
  wire [9:0] T_1304;
  wire  T_1306;
  wire [9:0] T_1312;
  wire [9:0] T_1313;
  wire  T_1315;
  wire [9:0] T_1321;
  wire [9:0] T_1322;
  wire  T_1324;
  wire [9:0] T_1330;
  wire [9:0] T_1331;
  wire  T_1333;
  wire [9:0] T_1339;
  wire [9:0] T_1340;
  wire  T_1342;
  wire  T_1350_0;
  wire  T_1350_1;
  wire  T_1350_2;
  wire  T_1350_3;
  wire  T_1350_4;
  wire  T_1350_5;
  wire  T_1350_6;
  wire  T_1350_7;
  wire  T_1350_8;
  wire  T_1350_9;
  wire  T_1350_10;
  wire  T_1350_11;
  wire  T_1350_12;
  wire  T_1350_13;
  wire  T_1350_14;
  wire  T_1350_15;
  wire  T_1350_16;
  wire  T_1350_17;
  wire  T_1350_18;
  wire  T_1350_19;
  wire  T_1350_20;
  wire  T_1350_21;
  wire  T_1350_22;
  wire  T_1350_23;
  wire  T_1350_24;
  wire  T_1350_25;
  wire  T_1355_0;
  wire  T_1355_1;
  wire  T_1355_2;
  wire  T_1355_3;
  wire  T_1355_4;
  wire  T_1355_5;
  wire  T_1355_6;
  wire  T_1355_7;
  wire  T_1355_8;
  wire  T_1355_9;
  wire  T_1355_10;
  wire  T_1355_11;
  wire  T_1355_12;
  wire  T_1355_13;
  wire  T_1355_14;
  wire  T_1355_15;
  wire  T_1355_16;
  wire  T_1355_17;
  wire  T_1355_18;
  wire  T_1355_19;
  wire  T_1355_20;
  wire  T_1355_21;
  wire  T_1355_22;
  wire  T_1355_23;
  wire  T_1355_24;
  wire  T_1355_25;
  wire  T_1360_0;
  wire  T_1360_1;
  wire  T_1360_2;
  wire  T_1360_3;
  wire  T_1360_4;
  wire  T_1360_5;
  wire  T_1360_6;
  wire  T_1360_7;
  wire  T_1360_8;
  wire  T_1360_9;
  wire  T_1360_10;
  wire  T_1360_11;
  wire  T_1360_12;
  wire  T_1360_13;
  wire  T_1360_14;
  wire  T_1360_15;
  wire  T_1360_16;
  wire  T_1360_17;
  wire  T_1360_18;
  wire  T_1360_19;
  wire  T_1360_20;
  wire  T_1360_21;
  wire  T_1360_22;
  wire  T_1360_23;
  wire  T_1360_24;
  wire  T_1360_25;
  wire  T_1365_0;
  wire  T_1365_1;
  wire  T_1365_2;
  wire  T_1365_3;
  wire  T_1365_4;
  wire  T_1365_5;
  wire  T_1365_6;
  wire  T_1365_7;
  wire  T_1365_8;
  wire  T_1365_9;
  wire  T_1365_10;
  wire  T_1365_11;
  wire  T_1365_12;
  wire  T_1365_13;
  wire  T_1365_14;
  wire  T_1365_15;
  wire  T_1365_16;
  wire  T_1365_17;
  wire  T_1365_18;
  wire  T_1365_19;
  wire  T_1365_20;
  wire  T_1365_21;
  wire  T_1365_22;
  wire  T_1365_23;
  wire  T_1365_24;
  wire  T_1365_25;
  wire  T_1370_0;
  wire  T_1370_1;
  wire  T_1370_2;
  wire  T_1370_3;
  wire  T_1370_4;
  wire  T_1370_5;
  wire  T_1370_6;
  wire  T_1370_7;
  wire  T_1370_8;
  wire  T_1370_9;
  wire  T_1370_10;
  wire  T_1370_11;
  wire  T_1370_12;
  wire  T_1370_13;
  wire  T_1370_14;
  wire  T_1370_15;
  wire  T_1370_16;
  wire  T_1370_17;
  wire  T_1370_18;
  wire  T_1370_19;
  wire  T_1370_20;
  wire  T_1370_21;
  wire  T_1370_22;
  wire  T_1370_23;
  wire  T_1370_24;
  wire  T_1370_25;
  wire  T_1375_0;
  wire  T_1375_1;
  wire  T_1375_2;
  wire  T_1375_3;
  wire  T_1375_4;
  wire  T_1375_5;
  wire  T_1375_6;
  wire  T_1375_7;
  wire  T_1375_8;
  wire  T_1375_9;
  wire  T_1375_10;
  wire  T_1375_11;
  wire  T_1375_12;
  wire  T_1375_13;
  wire  T_1375_14;
  wire  T_1375_15;
  wire  T_1375_16;
  wire  T_1375_17;
  wire  T_1375_18;
  wire  T_1375_19;
  wire  T_1375_20;
  wire  T_1375_21;
  wire  T_1375_22;
  wire  T_1375_23;
  wire  T_1375_24;
  wire  T_1375_25;
  wire  T_1380_0;
  wire  T_1380_1;
  wire  T_1380_2;
  wire  T_1380_3;
  wire  T_1380_4;
  wire  T_1380_5;
  wire  T_1380_6;
  wire  T_1380_7;
  wire  T_1380_8;
  wire  T_1380_9;
  wire  T_1380_10;
  wire  T_1380_11;
  wire  T_1380_12;
  wire  T_1380_13;
  wire  T_1380_14;
  wire  T_1380_15;
  wire  T_1380_16;
  wire  T_1380_17;
  wire  T_1380_18;
  wire  T_1380_19;
  wire  T_1380_20;
  wire  T_1380_21;
  wire  T_1380_22;
  wire  T_1380_23;
  wire  T_1380_24;
  wire  T_1380_25;
  wire  T_1385_0;
  wire  T_1385_1;
  wire  T_1385_2;
  wire  T_1385_3;
  wire  T_1385_4;
  wire  T_1385_5;
  wire  T_1385_6;
  wire  T_1385_7;
  wire  T_1385_8;
  wire  T_1385_9;
  wire  T_1385_10;
  wire  T_1385_11;
  wire  T_1385_12;
  wire  T_1385_13;
  wire  T_1385_14;
  wire  T_1385_15;
  wire  T_1385_16;
  wire  T_1385_17;
  wire  T_1385_18;
  wire  T_1385_19;
  wire  T_1385_20;
  wire  T_1385_21;
  wire  T_1385_22;
  wire  T_1385_23;
  wire  T_1385_24;
  wire  T_1385_25;
  wire  T_1547;
  wire  T_1548;
  wire  T_1549;
  wire  T_1550;
  wire [7:0] T_1554;
  wire [7:0] T_1558;
  wire [7:0] T_1562;
  wire [7:0] T_1566;
  wire [15:0] T_1567;
  wire [15:0] T_1568;
  wire [31:0] T_1569;
  wire [11:0] T_1593;
  wire [11:0] T_1597;
  wire  T_1599;
  wire  T_1612;
  wire [11:0] T_1613;
  wire [11:0] GEN_6;
  wire  T_1633;
  wire  T_1637;
  wire  T_1639;
  wire  T_1652;
  wire  T_1653;
  wire  GEN_7;
  wire [7:0] T_1673;
  wire  T_1675;
  wire [7:0] T_1677;
  wire  T_1679;
  wire  T_1692;
  wire [7:0] T_1693;
  wire [7:0] GEN_8;
  wire [7:0] T_1713;
  wire [7:0] T_1717;
  wire  T_1719;
  wire  T_1732;
  wire [7:0] T_1733;
  wire [7:0] GEN_9;
  wire [23:0] GEN_210;
  wire [23:0] T_1748;
  wire [23:0] GEN_211;
  wire [23:0] T_1752;
  wire [3:0] T_1753;
  wire [3:0] T_1757;
  wire  T_1759;
  wire  T_1772;
  wire [3:0] T_1773;
  wire [3:0] GEN_10;
  wire  T_1828;
  wire  T_1833;
  wire  T_1837;
  wire  T_1839;
  wire  T_1853;
  wire [1:0] GEN_212;
  wire [1:0] T_1868;
  wire [1:0] GEN_213;
  wire [1:0] T_1872;
  wire  T_1892;
  wire  GEN_11;
  wire  T_1932;
  wire  GEN_12;
  wire [1:0] GEN_214;
  wire [1:0] T_1948;
  wire [1:0] GEN_215;
  wire [1:0] T_1952;
  wire [1:0] T_1953;
  wire [1:0] T_1957;
  wire  T_1959;
  wire  T_1972;
  wire [1:0] T_1973;
  wire [1:0] GEN_13;
  wire  T_2012;
  wire  GEN_14;
  wire  T_2052;
  wire  GEN_15;
  wire [1:0] GEN_216;
  wire [1:0] T_2068;
  wire [1:0] GEN_217;
  wire [1:0] T_2072;
  wire  T_2092;
  wire [3:0] GEN_16;
  wire  T_2132;
  wire [31:0] GEN_218;
  wire [31:0] T_2228;
  wire  T_2252;
  wire [1:0] GEN_17;
  wire  T_2273;
  wire  T_2277;
  wire  T_2279;
  wire  T_2292;
  wire  T_2293;
  wire  GEN_18;
  wire [2:0] GEN_219;
  wire [2:0] T_2308;
  wire [2:0] GEN_220;
  wire [2:0] T_2312;
  wire  T_2313;
  wire  T_2317;
  wire  T_2319;
  wire  T_2332;
  wire  T_2333;
  wire  GEN_19;
  wire [3:0] GEN_221;
  wire [3:0] T_2348;
  wire [3:0] GEN_222;
  wire [3:0] T_2352;
  wire [3:0] T_2353;
  wire [3:0] T_2357;
  wire  T_2359;
  wire  T_2372;
  wire [3:0] T_2373;
  wire [3:0] GEN_20;
  wire [19:0] GEN_223;
  wire [19:0] T_2388;
  wire [19:0] GEN_224;
  wire [19:0] T_2392;
  wire  T_2412;
  wire [7:0] GEN_21;
  wire  T_2452;
  wire [7:0] GEN_22;
  wire [23:0] GEN_225;
  wire [23:0] T_2468;
  wire [23:0] GEN_226;
  wire [23:0] T_2472;
  wire  T_2488;
  wire [7:0] T_2508;
  wire [30:0] T_2552;
  wire [31:0] GEN_227;
  wire [31:0] T_2588;
  wire [31:0] GEN_228;
  wire [31:0] T_2592;
  wire  T_2612;
  wire  GEN_23;
  wire  T_2634;
  wire  T_2636;
  wire  T_2638;
  wire  T_2639;
  wire  T_2641;
  wire  T_2649;
  wire  T_2651;
  wire  T_2653;
  wire  T_2655;
  wire  T_2657;
  wire  T_2659;
  wire  T_2670;
  wire  T_2671;
  wire  T_2673;
  wire  T_2675;
  wire  T_2676;
  wire  T_2678;
  wire  T_2692;
  wire  T_2693;
  wire  T_2694;
  wire  T_2695;
  wire  T_2697;
  wire  T_2702;
  wire  T_2703;
  wire  T_2704;
  wire  T_2706;
  wire  T_2708;
  wire  T_2709;
  wire  T_2710;
  wire  T_2712;
  wire  T_2714;
  wire  T_2716;
  wire  T_2718;
  wire  T_2720;
  wire  T_2740;
  wire  T_2741;
  wire  T_2743;
  wire  T_2745;
  wire  T_2746;
  wire  T_2748;
  wire  T_2790_0;
  wire  T_2790_1;
  wire  T_2790_2;
  wire  T_2790_3;
  wire  T_2790_4;
  wire  T_2790_5;
  wire  T_2790_6;
  wire  T_2790_7;
  wire  T_2790_8;
  wire  T_2790_9;
  wire  T_2790_10;
  wire  T_2790_11;
  wire  T_2790_12;
  wire  T_2790_13;
  wire  T_2790_14;
  wire  T_2790_15;
  wire  T_2790_16;
  wire  T_2790_17;
  wire  T_2790_18;
  wire  T_2790_19;
  wire  T_2790_20;
  wire  T_2790_21;
  wire  T_2790_22;
  wire  T_2790_23;
  wire  T_2790_24;
  wire  T_2790_25;
  wire  T_2790_26;
  wire  T_2790_27;
  wire  T_2790_28;
  wire  T_2790_29;
  wire  T_2790_30;
  wire  T_2790_31;
  wire  T_2828;
  wire  T_2831;
  wire  T_2833;
  wire  T_2843;
  wire  T_2847;
  wire  T_2851;
  wire  T_2863;
  wire  T_2865;
  wire  T_2868;
  wire  T_2870;
  wire  T_2885;
  wire  T_2886;
  wire  T_2887;
  wire  T_2889;
  wire  T_2895;
  wire  T_2896;
  wire  T_2898;
  wire  T_2901;
  wire  T_2902;
  wire  T_2904;
  wire  T_2908;
  wire  T_2912;
  wire  T_2933;
  wire  T_2935;
  wire  T_2938;
  wire  T_2940;
  wire  T_2982_0;
  wire  T_2982_1;
  wire  T_2982_2;
  wire  T_2982_3;
  wire  T_2982_4;
  wire  T_2982_5;
  wire  T_2982_6;
  wire  T_2982_7;
  wire  T_2982_8;
  wire  T_2982_9;
  wire  T_2982_10;
  wire  T_2982_11;
  wire  T_2982_12;
  wire  T_2982_13;
  wire  T_2982_14;
  wire  T_2982_15;
  wire  T_2982_16;
  wire  T_2982_17;
  wire  T_2982_18;
  wire  T_2982_19;
  wire  T_2982_20;
  wire  T_2982_21;
  wire  T_2982_22;
  wire  T_2982_23;
  wire  T_2982_24;
  wire  T_2982_25;
  wire  T_2982_26;
  wire  T_2982_27;
  wire  T_2982_28;
  wire  T_2982_29;
  wire  T_2982_30;
  wire  T_2982_31;
  wire  T_3020;
  wire  T_3023;
  wire  T_3025;
  wire  T_3035;
  wire  T_3039;
  wire  T_3043;
  wire  T_3055;
  wire  T_3057;
  wire  T_3060;
  wire  T_3062;
  wire  T_3077;
  wire  T_3078;
  wire  T_3079;
  wire  T_3081;
  wire  T_3087;
  wire  T_3088;
  wire  T_3090;
  wire  T_3093;
  wire  T_3094;
  wire  T_3096;
  wire  T_3100;
  wire  T_3104;
  wire  T_3125;
  wire  T_3127;
  wire  T_3130;
  wire  T_3132;
  wire  T_3174_0;
  wire  T_3174_1;
  wire  T_3174_2;
  wire  T_3174_3;
  wire  T_3174_4;
  wire  T_3174_5;
  wire  T_3174_6;
  wire  T_3174_7;
  wire  T_3174_8;
  wire  T_3174_9;
  wire  T_3174_10;
  wire  T_3174_11;
  wire  T_3174_12;
  wire  T_3174_13;
  wire  T_3174_14;
  wire  T_3174_15;
  wire  T_3174_16;
  wire  T_3174_17;
  wire  T_3174_18;
  wire  T_3174_19;
  wire  T_3174_20;
  wire  T_3174_21;
  wire  T_3174_22;
  wire  T_3174_23;
  wire  T_3174_24;
  wire  T_3174_25;
  wire  T_3174_26;
  wire  T_3174_27;
  wire  T_3174_28;
  wire  T_3174_29;
  wire  T_3174_30;
  wire  T_3174_31;
  wire  T_3212;
  wire  T_3215;
  wire  T_3217;
  wire  T_3227;
  wire  T_3231;
  wire  T_3235;
  wire  T_3247;
  wire  T_3249;
  wire  T_3252;
  wire  T_3254;
  wire  T_3269;
  wire  T_3270;
  wire  T_3271;
  wire  T_3273;
  wire  T_3279;
  wire  T_3280;
  wire  T_3282;
  wire  T_3285;
  wire  T_3286;
  wire  T_3288;
  wire  T_3292;
  wire  T_3296;
  wire  T_3317;
  wire  T_3319;
  wire  T_3322;
  wire  T_3324;
  wire  T_3366_0;
  wire  T_3366_1;
  wire  T_3366_2;
  wire  T_3366_3;
  wire  T_3366_4;
  wire  T_3366_5;
  wire  T_3366_6;
  wire  T_3366_7;
  wire  T_3366_8;
  wire  T_3366_9;
  wire  T_3366_10;
  wire  T_3366_11;
  wire  T_3366_12;
  wire  T_3366_13;
  wire  T_3366_14;
  wire  T_3366_15;
  wire  T_3366_16;
  wire  T_3366_17;
  wire  T_3366_18;
  wire  T_3366_19;
  wire  T_3366_20;
  wire  T_3366_21;
  wire  T_3366_22;
  wire  T_3366_23;
  wire  T_3366_24;
  wire  T_3366_25;
  wire  T_3366_26;
  wire  T_3366_27;
  wire  T_3366_28;
  wire  T_3366_29;
  wire  T_3366_30;
  wire  T_3366_31;
  wire  T_3401;
  wire  T_3402;
  wire  T_3403;
  wire  T_3404;
  wire  T_3405;
  wire [1:0] T_3411;
  wire [1:0] T_3412;
  wire [2:0] T_3413;
  wire [4:0] T_3414;
  wire  GEN_0;
  wire  GEN_24;
  wire  GEN_25;
  wire  GEN_26;
  wire  GEN_27;
  wire  GEN_28;
  wire  GEN_29;
  wire  GEN_30;
  wire  GEN_31;
  wire  GEN_32;
  wire  GEN_33;
  wire  GEN_34;
  wire  GEN_35;
  wire  GEN_36;
  wire  GEN_37;
  wire  GEN_38;
  wire  GEN_39;
  wire  GEN_40;
  wire  GEN_41;
  wire  GEN_42;
  wire  GEN_43;
  wire  GEN_44;
  wire  GEN_45;
  wire  GEN_46;
  wire  GEN_47;
  wire  GEN_48;
  wire  GEN_49;
  wire  GEN_50;
  wire  GEN_51;
  wire  GEN_52;
  wire  GEN_53;
  wire  GEN_54;
  wire  GEN_1;
  wire  GEN_55;
  wire  GEN_56;
  wire  GEN_57;
  wire  GEN_58;
  wire  GEN_59;
  wire  GEN_60;
  wire  GEN_61;
  wire  GEN_62;
  wire  GEN_63;
  wire  GEN_64;
  wire  GEN_65;
  wire  GEN_66;
  wire  GEN_67;
  wire  GEN_68;
  wire  GEN_69;
  wire  GEN_70;
  wire  GEN_71;
  wire  GEN_72;
  wire  GEN_73;
  wire  GEN_74;
  wire  GEN_75;
  wire  GEN_76;
  wire  GEN_77;
  wire  GEN_78;
  wire  GEN_79;
  wire  GEN_80;
  wire  GEN_81;
  wire  GEN_82;
  wire  GEN_83;
  wire  GEN_84;
  wire  GEN_85;
  wire  T_3431;
  wire  GEN_2;
  wire  GEN_86;
  wire  GEN_87;
  wire  GEN_88;
  wire  GEN_89;
  wire  GEN_90;
  wire  GEN_91;
  wire  GEN_92;
  wire  GEN_93;
  wire  GEN_94;
  wire  GEN_95;
  wire  GEN_96;
  wire  GEN_97;
  wire  GEN_98;
  wire  GEN_99;
  wire  GEN_100;
  wire  GEN_101;
  wire  GEN_102;
  wire  GEN_103;
  wire  GEN_104;
  wire  GEN_105;
  wire  GEN_106;
  wire  GEN_107;
  wire  GEN_108;
  wire  GEN_109;
  wire  GEN_110;
  wire  GEN_111;
  wire  GEN_112;
  wire  GEN_113;
  wire  GEN_114;
  wire  GEN_115;
  wire  GEN_116;
  wire  GEN_3;
  wire  GEN_117;
  wire  GEN_118;
  wire  GEN_119;
  wire  GEN_120;
  wire  GEN_121;
  wire  GEN_122;
  wire  GEN_123;
  wire  GEN_124;
  wire  GEN_125;
  wire  GEN_126;
  wire  GEN_127;
  wire  GEN_128;
  wire  GEN_129;
  wire  GEN_130;
  wire  GEN_131;
  wire  GEN_132;
  wire  GEN_133;
  wire  GEN_134;
  wire  GEN_135;
  wire  GEN_136;
  wire  GEN_137;
  wire  GEN_138;
  wire  GEN_139;
  wire  GEN_140;
  wire  GEN_141;
  wire  GEN_142;
  wire  GEN_143;
  wire  GEN_144;
  wire  GEN_145;
  wire  GEN_146;
  wire  GEN_147;
  wire  T_3434;
  wire  T_3435;
  wire  T_3436;
  wire  T_3437;
  wire  T_3438;
  wire [31:0] T_3440;
  wire [1:0] T_3441;
  wire [3:0] T_3443;
  wire [1:0] T_3444;
  wire [1:0] T_3445;
  wire [3:0] T_3446;
  wire [7:0] T_3447;
  wire [1:0] T_3449;
  wire [3:0] T_3450;
  wire [7:0] T_3454;
  wire [15:0] T_3455;
  wire [1:0] T_3456;
  wire [1:0] T_3457;
  wire [3:0] T_3458;
  wire [1:0] T_3459;
  wire [3:0] T_3461;
  wire [7:0] T_3462;
  wire [1:0] T_3466;
  wire [3:0] T_3468;
  wire [7:0] T_3469;
  wire [15:0] T_3470;
  wire [31:0] T_3471;
  wire [31:0] T_3472;
  wire  T_3507;
  wire  T_3508;
  wire  T_3509;
  wire  T_3510;
  wire  T_3513;
  wire  T_3514;
  wire  T_3516;
  wire  T_3517;
  wire  T_3518;
  wire  T_3520;
  wire  T_3524;
  wire  T_3526;
  wire  T_3529;
  wire  T_3530;
  wire  T_3536;
  wire  T_3540;
  wire  T_3546;
  wire  T_3589;
  wire  T_3590;
  wire  T_3596;
  wire  T_3600;
  wire  T_3606;
  wire  T_3609;
  wire  T_3610;
  wire  T_3616;
  wire  T_3620;
  wire  T_3626;
  wire  T_3629;
  wire  T_3630;
  wire  T_3636;
  wire  T_3640;
  wire  T_3646;
  wire  T_3709;
  wire  T_3710;
  wire  T_3716;
  wire  T_3720;
  wire  T_3726;
  wire  T_3729;
  wire  T_3730;
  wire  T_3736;
  wire  T_3740;
  wire  T_3746;
  wire  T_3829;
  wire  T_3830;
  wire  T_3836;
  wire  T_3840;
  wire  T_3846;
  wire  T_3869;
  wire  T_3870;
  wire  T_3876;
  wire  T_3880;
  wire  T_3886;
  wire  T_3889;
  wire  T_3890;
  wire  T_3896;
  wire  T_3900;
  wire  T_3906;
  wire  T_3909;
  wire  T_3910;
  wire  T_3916;
  wire  T_3920;
  wire  T_3926;
  wire  T_3929;
  wire  T_3930;
  wire  T_3936;
  wire  T_3940;
  wire  T_3946;
  wire  T_4069;
  wire  T_4070;
  wire  T_4076;
  wire  T_4080;
  wire  T_4086;
  wire  T_4089;
  wire  T_4090;
  wire  T_4096;
  wire  T_4100;
  wire  T_4106;
  wire  T_4155;
  wire  T_4157;
  wire  T_4159;
  wire  T_4161;
  wire  T_4163;
  wire  T_4165;
  wire  T_4167;
  wire  T_4169;
  wire  T_4175;
  wire  T_4177;
  wire  T_4179;
  wire  T_4181;
  wire  T_4183;
  wire  T_4185;
  wire  T_4187;
  wire  T_4189;
  wire  T_4191;
  wire  T_4193;
  wire  T_4195;
  wire  T_4197;
  wire  T_4199;
  wire  T_4201;
  wire  T_4203;
  wire  T_4205;
  wire  T_4211;
  wire  T_4213;
  wire  T_4215;
  wire  T_4217;
  wire  T_4219;
  wire  T_4221;
  wire  T_4223;
  wire  T_4225;
  wire  T_4231;
  wire  T_4232;
  wire  T_4234;
  wire  T_4235;
  wire  T_4237;
  wire  T_4238;
  wire  T_4240;
  wire  T_4241;
  wire  T_4244;
  wire  T_4247;
  wire  T_4250;
  wire  T_4253;
  wire  T_4255;
  wire  T_4256;
  wire  T_4258;
  wire  T_4259;
  wire  T_4261;
  wire  T_4262;
  wire  T_4264;
  wire  T_4265;
  wire  T_4267;
  wire  T_4268;
  wire  T_4269;
  wire  T_4271;
  wire  T_4272;
  wire  T_4273;
  wire  T_4275;
  wire  T_4276;
  wire  T_4277;
  wire  T_4279;
  wire  T_4280;
  wire  T_4281;
  wire  T_4285;
  wire  T_4289;
  wire  T_4293;
  wire  T_4297;
  wire  T_4300;
  wire  T_4301;
  wire  T_4304;
  wire  T_4305;
  wire  T_4308;
  wire  T_4309;
  wire  T_4312;
  wire  T_4313;
  wire  T_4315;
  wire  T_4316;
  wire  T_4317;
  wire  T_4319;
  wire  T_4320;
  wire  T_4321;
  wire  T_4323;
  wire  T_4324;
  wire  T_4325;
  wire  T_4327;
  wire  T_4328;
  wire  T_4329;
  wire  T_4331;
  wire  T_4333;
  wire  T_4335;
  wire  T_4337;
  wire  T_4339;
  wire  T_4341;
  wire  T_4343;
  wire  T_4345;
  wire  T_4347;
  wire  T_4348;
  wire  T_4350;
  wire  T_4351;
  wire  T_4353;
  wire  T_4354;
  wire  T_4356;
  wire  T_4357;
  wire  T_4360;
  wire  T_4363;
  wire  T_4366;
  wire  T_4369;
  wire  T_4371;
  wire  T_4372;
  wire  T_4374;
  wire  T_4375;
  wire  T_4377;
  wire  T_4378;
  wire  T_4380;
  wire  T_4381;
  wire  T_4422_0;
  wire  T_4422_1;
  wire  T_4422_2;
  wire  T_4422_3;
  wire  T_4422_4;
  wire  T_4422_5;
  wire  T_4422_6;
  wire  T_4422_7;
  wire  T_4422_8;
  wire  T_4422_9;
  wire  T_4422_10;
  wire  T_4422_11;
  wire  T_4422_12;
  wire  T_4422_13;
  wire  T_4422_14;
  wire  T_4422_15;
  wire  T_4422_16;
  wire  T_4422_17;
  wire  T_4422_18;
  wire  T_4422_19;
  wire  T_4422_20;
  wire  T_4422_21;
  wire  T_4422_22;
  wire  T_4422_23;
  wire  T_4422_24;
  wire  T_4422_25;
  wire  T_4422_26;
  wire  T_4422_27;
  wire  T_4422_28;
  wire  T_4422_29;
  wire  T_4422_30;
  wire  T_4422_31;
  wire [31:0] T_4493_0;
  wire [31:0] T_4493_1;
  wire [31:0] T_4493_2;
  wire [31:0] T_4493_3;
  wire [31:0] T_4493_4;
  wire [31:0] T_4493_5;
  wire [31:0] T_4493_6;
  wire [31:0] T_4493_7;
  wire [31:0] T_4493_8;
  wire [31:0] T_4493_9;
  wire [31:0] T_4493_10;
  wire [31:0] T_4493_11;
  wire [31:0] T_4493_12;
  wire [31:0] T_4493_13;
  wire [31:0] T_4493_14;
  wire [31:0] T_4493_15;
  wire [31:0] T_4493_16;
  wire [31:0] T_4493_17;
  wire [31:0] T_4493_18;
  wire [31:0] T_4493_19;
  wire [31:0] T_4493_20;
  wire [31:0] T_4493_21;
  wire [31:0] T_4493_22;
  wire [31:0] T_4493_23;
  wire [31:0] T_4493_24;
  wire [31:0] T_4493_25;
  wire [31:0] T_4493_26;
  wire [31:0] T_4493_27;
  wire [31:0] T_4493_28;
  wire [31:0] T_4493_29;
  wire [31:0] T_4493_30;
  wire [31:0] T_4493_31;
  wire  GEN_4;
  wire  GEN_148;
  wire  GEN_149;
  wire  GEN_150;
  wire  GEN_151;
  wire  GEN_152;
  wire  GEN_153;
  wire  GEN_154;
  wire  GEN_155;
  wire  GEN_156;
  wire  GEN_157;
  wire  GEN_158;
  wire  GEN_159;
  wire  GEN_160;
  wire  GEN_161;
  wire  GEN_162;
  wire  GEN_163;
  wire  GEN_164;
  wire  GEN_165;
  wire  GEN_166;
  wire  GEN_167;
  wire  GEN_168;
  wire  GEN_169;
  wire  GEN_170;
  wire  GEN_171;
  wire  GEN_172;
  wire  GEN_173;
  wire  GEN_174;
  wire  GEN_175;
  wire  GEN_176;
  wire  GEN_177;
  wire  GEN_178;
  wire [31:0] GEN_5;
  wire [31:0] GEN_179;
  wire [31:0] GEN_180;
  wire [31:0] GEN_181;
  wire [31:0] GEN_182;
  wire [31:0] GEN_183;
  wire [31:0] GEN_184;
  wire [31:0] GEN_185;
  wire [31:0] GEN_186;
  wire [31:0] GEN_187;
  wire [31:0] GEN_188;
  wire [31:0] GEN_189;
  wire [31:0] GEN_190;
  wire [31:0] GEN_191;
  wire [31:0] GEN_192;
  wire [31:0] GEN_193;
  wire [31:0] GEN_194;
  wire [31:0] GEN_195;
  wire [31:0] GEN_196;
  wire [31:0] GEN_197;
  wire [31:0] GEN_198;
  wire [31:0] GEN_199;
  wire [31:0] GEN_200;
  wire [31:0] GEN_201;
  wire [31:0] GEN_202;
  wire [31:0] GEN_203;
  wire [31:0] GEN_204;
  wire [31:0] GEN_205;
  wire [31:0] GEN_206;
  wire [31:0] GEN_207;
  wire [31:0] GEN_208;
  wire [31:0] GEN_209;
  wire [31:0] T_4530;
  wire [1:0] T_4531;
  wire [4:0] T_4533;
  wire [2:0] T_4534;
  wire [2:0] T_4545_opcode;
  wire [1:0] T_4545_param;
  wire [2:0] T_4545_size;
  wire [4:0] T_4545_source;
  wire  T_4545_sink;
  wire [1:0] T_4545_addr_lo;
  wire [31:0] T_4545_data;
  wire  T_4545_error;
  wire [2:0] GEN_229 = 3'b0;
  reg [31:0] GEN_254;
  wire [1:0] GEN_230 = 2'b0;
  reg [31:0] GEN_255;
  wire [2:0] GEN_231 = 3'b0;
  reg [31:0] GEN_256;
  wire [4:0] GEN_232 = 5'b0;
  reg [31:0] GEN_257;
  wire [28:0] GEN_233 = 29'b0;
  reg [31:0] GEN_258;
  wire [3:0] GEN_234 = 4'b0;
  reg [31:0] GEN_259;
  wire [31:0] GEN_235 = 32'b0;
  reg [31:0] GEN_260;
  sirv_qspi_fifo fifo (
    .clock(fifo_clock),
    .reset(fifo_reset),
    .io_ctrl_fmt_proto(fifo_io_ctrl_fmt_proto),
    .io_ctrl_fmt_endian(fifo_io_ctrl_fmt_endian),
    .io_ctrl_fmt_iodir(fifo_io_ctrl_fmt_iodir),
    .io_ctrl_fmt_len(fifo_io_ctrl_fmt_len),
    .io_ctrl_cs_mode(fifo_io_ctrl_cs_mode),
    .io_ctrl_wm_tx(fifo_io_ctrl_wm_tx),
    .io_ctrl_wm_rx(fifo_io_ctrl_wm_rx),
    .io_link_tx_ready(fifo_io_link_tx_ready),
    .io_link_tx_valid(fifo_io_link_tx_valid),
    .io_link_tx_bits(fifo_io_link_tx_bits),
    .io_link_rx_valid(fifo_io_link_rx_valid),
    .io_link_rx_bits(fifo_io_link_rx_bits),
    .io_link_cnt(fifo_io_link_cnt),
    .io_link_fmt_proto(fifo_io_link_fmt_proto),
    .io_link_fmt_endian(fifo_io_link_fmt_endian),
    .io_link_fmt_iodir(fifo_io_link_fmt_iodir),
    .io_link_cs_set(fifo_io_link_cs_set),
    .io_link_cs_clear(fifo_io_link_cs_clear),
    .io_link_cs_hold(fifo_io_link_cs_hold),
    .io_link_active(fifo_io_link_active),
    .io_link_lock(fifo_io_link_lock),
    .io_tx_ready(fifo_io_tx_ready),
    .io_tx_valid(fifo_io_tx_valid),
    .io_tx_bits(fifo_io_tx_bits),
    .io_rx_ready(fifo_io_rx_ready),
    .io_rx_valid(fifo_io_rx_valid),
    .io_rx_bits(fifo_io_rx_bits),
    .io_ip_txwm(fifo_io_ip_txwm),
    .io_ip_rxwm(fifo_io_ip_rxwm)
  );
  sirv_qspi_media_2 mac (
    .clock(mac_clock),
    .reset(mac_reset),
    .io_port_sck(mac_io_port_sck),
    .io_port_dq_0_i(mac_io_port_dq_0_i),
    .io_port_dq_0_o(mac_io_port_dq_0_o),
    .io_port_dq_0_oe(mac_io_port_dq_0_oe),
    .io_port_dq_1_i(mac_io_port_dq_1_i),
    .io_port_dq_1_o(mac_io_port_dq_1_o),
    .io_port_dq_1_oe(mac_io_port_dq_1_oe),
    .io_port_dq_2_i(mac_io_port_dq_2_i),
    .io_port_dq_2_o(mac_io_port_dq_2_o),
    .io_port_dq_2_oe(mac_io_port_dq_2_oe),
    .io_port_dq_3_i(mac_io_port_dq_3_i),
    .io_port_dq_3_o(mac_io_port_dq_3_o),
    .io_port_dq_3_oe(mac_io_port_dq_3_oe),
    .io_port_cs_0(mac_io_port_cs_0),
    .io_ctrl_sck_div(mac_io_ctrl_sck_div),
    .io_ctrl_sck_pol(mac_io_ctrl_sck_pol),
    .io_ctrl_sck_pha(mac_io_ctrl_sck_pha),
    .io_ctrl_dla_cssck(mac_io_ctrl_dla_cssck),
    .io_ctrl_dla_sckcs(mac_io_ctrl_dla_sckcs),
    .io_ctrl_dla_intercs(mac_io_ctrl_dla_intercs),
    .io_ctrl_dla_interxfr(mac_io_ctrl_dla_interxfr),
    .io_ctrl_cs_id(mac_io_ctrl_cs_id),
    .io_ctrl_cs_dflt_0(mac_io_ctrl_cs_dflt_0),
    .io_link_tx_ready(mac_io_link_tx_ready),
    .io_link_tx_valid(mac_io_link_tx_valid),
    .io_link_tx_bits(mac_io_link_tx_bits),
    .io_link_rx_valid(mac_io_link_rx_valid),
    .io_link_rx_bits(mac_io_link_rx_bits),
    .io_link_cnt(mac_io_link_cnt),
    .io_link_fmt_proto(mac_io_link_fmt_proto),
    .io_link_fmt_endian(mac_io_link_fmt_endian),
    .io_link_fmt_iodir(mac_io_link_fmt_iodir),
    .io_link_cs_set(mac_io_link_cs_set),
    .io_link_cs_clear(mac_io_link_cs_clear),
    .io_link_cs_hold(mac_io_link_cs_hold),
    .io_link_active(mac_io_link_active)
  );
  assign io_port_sck = mac_io_port_sck;
  assign io_port_dq_0_o = mac_io_port_dq_0_o;
  assign io_port_dq_0_oe = mac_io_port_dq_0_oe;
  assign io_port_dq_1_o = mac_io_port_dq_1_o;
  assign io_port_dq_1_oe = mac_io_port_dq_1_oe;
  assign io_port_dq_2_o = mac_io_port_dq_2_o;
  assign io_port_dq_2_oe = mac_io_port_dq_2_oe;
  assign io_port_dq_3_o = mac_io_port_dq_3_o;
  assign io_port_dq_3_oe = mac_io_port_dq_3_oe;
  assign io_port_cs_0 = mac_io_port_cs_0;
  assign io_tl_i_0_0 = T_1032;
  assign io_tl_r_0_a_ready = T_1063_ready;
  assign io_tl_r_0_b_valid = 1'h0;
  assign io_tl_r_0_b_bits_opcode = GEN_229;
  assign io_tl_r_0_b_bits_param = GEN_230;
  assign io_tl_r_0_b_bits_size = GEN_231;
  assign io_tl_r_0_b_bits_source = GEN_232;
  assign io_tl_r_0_b_bits_address = GEN_233;
  assign io_tl_r_0_b_bits_mask = GEN_234;
  assign io_tl_r_0_b_bits_data = GEN_235;
  assign io_tl_r_0_c_ready = 1'h1;
  assign io_tl_r_0_d_valid = T_1102_valid;
  assign io_tl_r_0_d_bits_opcode = {{2'd0}, T_1102_bits_read};
  assign io_tl_r_0_d_bits_param = T_4545_param;
  assign io_tl_r_0_d_bits_size = T_4545_size;
  assign io_tl_r_0_d_bits_source = T_4545_source;
  assign io_tl_r_0_d_bits_sink = T_4545_sink;
  assign io_tl_r_0_d_bits_addr_lo = T_4545_addr_lo;
  assign io_tl_r_0_d_bits_data = T_1102_bits_data;
  assign io_tl_r_0_d_bits_error = T_4545_error;
  assign io_tl_r_0_e_ready = 1'h1;
  assign T_955_fmt_proto = 2'h0;
  assign T_955_fmt_endian = 1'h0;
  assign T_955_fmt_iodir = 1'h0;
  assign T_955_fmt_len = 4'h8;
  assign T_955_sck_div = 12'h3;
  assign T_955_sck_pol = 1'h0;
  assign T_955_sck_pha = 1'h0;
  assign T_955_cs_id = 1'h0;
  assign T_955_cs_dflt_0 = 1'h1;
  assign T_955_cs_mode = 2'h0;
  assign T_955_dla_cssck = 8'h1;
  assign T_955_dla_sckcs = 8'h1;
  assign T_955_dla_intercs = 8'h1;
  assign T_955_dla_interxfr = 8'h0;
  assign T_955_wm_tx = 4'h0;
  assign T_955_wm_rx = 4'h0;
  assign fifo_clock = clock;
  assign fifo_reset = reset;
  assign fifo_io_ctrl_fmt_proto = ctrl_fmt_proto;
  assign fifo_io_ctrl_fmt_endian = ctrl_fmt_endian;
  assign fifo_io_ctrl_fmt_iodir = ctrl_fmt_iodir;
  assign fifo_io_ctrl_fmt_len = ctrl_fmt_len;
  assign fifo_io_ctrl_cs_mode = ctrl_cs_mode;
  assign fifo_io_ctrl_wm_tx = ctrl_wm_tx;
  assign fifo_io_ctrl_wm_rx = ctrl_wm_rx;
  assign fifo_io_link_tx_ready = mac_io_link_tx_ready;
  assign fifo_io_link_rx_valid = mac_io_link_rx_valid;
  assign fifo_io_link_rx_bits = mac_io_link_rx_bits;
  assign fifo_io_link_active = mac_io_link_active;
  assign fifo_io_tx_valid = T_2132;
  assign fifo_io_tx_bits = T_1693;
  assign fifo_io_rx_ready = T_2488;
  assign mac_clock = clock;
  assign mac_reset = reset;
  assign mac_io_port_dq_0_i = io_port_dq_0_i;
  assign mac_io_port_dq_1_i = io_port_dq_1_i;
  assign mac_io_port_dq_2_i = io_port_dq_2_i;
  assign mac_io_port_dq_3_i = io_port_dq_3_i;
  assign mac_io_ctrl_sck_div = ctrl_sck_div;
  assign mac_io_ctrl_sck_pol = ctrl_sck_pol;
  assign mac_io_ctrl_sck_pha = ctrl_sck_pha;
  assign mac_io_ctrl_dla_cssck = ctrl_dla_cssck;
  assign mac_io_ctrl_dla_sckcs = ctrl_dla_sckcs;
  assign mac_io_ctrl_dla_intercs = ctrl_dla_intercs;
  assign mac_io_ctrl_dla_interxfr = ctrl_dla_interxfr;
  assign mac_io_ctrl_cs_id = ctrl_cs_id;
  assign mac_io_ctrl_cs_dflt_0 = ctrl_cs_dflt_0;
  assign mac_io_link_tx_valid = fifo_io_link_tx_valid;
  assign mac_io_link_tx_bits = fifo_io_link_tx_bits;
  assign mac_io_link_cnt = fifo_io_link_cnt;
  assign mac_io_link_fmt_proto = fifo_io_link_fmt_proto;
  assign mac_io_link_fmt_endian = fifo_io_link_fmt_endian;
  assign mac_io_link_fmt_iodir = fifo_io_link_fmt_iodir;
  assign mac_io_link_cs_set = fifo_io_link_cs_set;
  assign mac_io_link_cs_clear = fifo_io_link_cs_clear;
  assign mac_io_link_cs_hold = fifo_io_link_cs_hold;
  assign T_1021_txwm = T_1027;
  assign T_1021_rxwm = T_1026;
  assign T_1025 = 2'h0;
  assign T_1026 = T_1025[0];
  assign T_1027 = T_1025[1];
  assign T_1030 = fifo_io_ip_txwm & ie_txwm;
  assign T_1031 = fifo_io_ip_rxwm & ie_rxwm;
  assign T_1032 = T_1030 | T_1031;
  assign T_1036 = fifo_io_tx_ready == 1'h0;
  assign T_1039 = fifo_io_rx_valid == 1'h0;
  assign T_1063_ready = T_3435;
  assign T_1063_valid = io_tl_r_0_a_valid;
  assign T_1063_bits_read = T_1080;
  assign T_1063_bits_index = T_1081[9:0];
  assign T_1063_bits_data = io_tl_r_0_a_bits_data;
  assign T_1063_bits_mask = io_tl_r_0_a_bits_mask;
  assign T_1063_bits_extra = T_1084;
  assign T_1080 = io_tl_r_0_a_bits_opcode == 3'h4;
  assign T_1081 = io_tl_r_0_a_bits_address[28:2];
  assign T_1082 = io_tl_r_0_a_bits_address[1:0];
  assign T_1083 = {T_1082,io_tl_r_0_a_bits_source};
  assign T_1084 = {T_1083,io_tl_r_0_a_bits_size};
  assign T_1102_ready = io_tl_r_0_d_ready;
  assign T_1102_valid = T_3438;
  assign T_1102_bits_read = T_1138_bits_read;
  assign T_1102_bits_data = T_4530;
  assign T_1102_bits_extra = T_1138_bits_extra;
  assign T_1138_ready = T_3437;
  assign T_1138_valid = T_3436;
  assign T_1138_bits_read = T_1063_bits_read;
  assign T_1138_bits_index = T_1063_bits_index;
  assign T_1138_bits_data = T_1063_bits_data;
  assign T_1138_bits_mask = T_1063_bits_mask;
  assign T_1138_bits_extra = T_1063_bits_extra;
  assign T_1223 = T_1138_bits_index & 10'h3e0;
  assign T_1225 = T_1223 == 10'h0;
  assign T_1231 = T_1138_bits_index ^ 10'h5;
  assign T_1232 = T_1231 & 10'h3e0;
  assign T_1234 = T_1232 == 10'h0;
  assign T_1240 = T_1138_bits_index ^ 10'ha;
  assign T_1241 = T_1240 & 10'h3e0;
  assign T_1243 = T_1241 == 10'h0;
  assign T_1249 = T_1138_bits_index ^ 10'h14;
  assign T_1250 = T_1249 & 10'h3e0;
  assign T_1252 = T_1250 == 10'h0;
  assign T_1258 = T_1138_bits_index ^ 10'h1d;
  assign T_1259 = T_1258 & 10'h3e0;
  assign T_1261 = T_1259 == 10'h0;
  assign T_1267 = T_1138_bits_index ^ 10'h1;
  assign T_1268 = T_1267 & 10'h3e0;
  assign T_1270 = T_1268 == 10'h0;
  assign T_1276 = T_1138_bits_index ^ 10'h6;
  assign T_1277 = T_1276 & 10'h3e0;
  assign T_1279 = T_1277 == 10'h0;
  assign T_1285 = T_1138_bits_index ^ 10'h1c;
  assign T_1286 = T_1285 & 10'h3e0;
  assign T_1288 = T_1286 == 10'h0;
  assign T_1294 = T_1138_bits_index ^ 10'h15;
  assign T_1295 = T_1294 & 10'h3e0;
  assign T_1297 = T_1295 == 10'h0;
  assign T_1303 = T_1138_bits_index ^ 10'h12;
  assign T_1304 = T_1303 & 10'h3e0;
  assign T_1306 = T_1304 == 10'h0;
  assign T_1312 = T_1138_bits_index ^ 10'h10;
  assign T_1313 = T_1312 & 10'h3e0;
  assign T_1315 = T_1313 == 10'h0;
  assign T_1321 = T_1138_bits_index ^ 10'hb;
  assign T_1322 = T_1321 & 10'h3e0;
  assign T_1324 = T_1322 == 10'h0;
  assign T_1330 = T_1138_bits_index ^ 10'h13;
  assign T_1331 = T_1330 & 10'h3e0;
  assign T_1333 = T_1331 == 10'h0;
  assign T_1339 = T_1138_bits_index ^ 10'h4;
  assign T_1340 = T_1339 & 10'h3e0;
  assign T_1342 = T_1340 == 10'h0;
  assign T_1350_0 = T_3510;
  assign T_1350_1 = T_3610;
  assign T_1350_2 = T_4155;
  assign T_1350_3 = T_4163;
  assign T_1350_4 = T_3910;
  assign T_1350_5 = T_4175;
  assign T_1350_6 = T_4183;
  assign T_1350_7 = T_4191;
  assign T_1350_8 = T_4199;
  assign T_1350_9 = T_3630;
  assign T_1350_10 = T_4211;
  assign T_1350_11 = T_4219;
  assign T_1350_12 = T_3930;
  assign T_1350_13 = T_4232;
  assign T_1350_14 = T_4244;
  assign T_1350_15 = T_4256;
  assign T_1350_16 = T_4269;
  assign T_1350_17 = T_4285;
  assign T_1350_18 = T_4301;
  assign T_1350_19 = T_4317;
  assign T_1350_20 = T_4331;
  assign T_1350_21 = T_4339;
  assign T_1350_22 = T_4348;
  assign T_1350_23 = T_4360;
  assign T_1350_24 = T_4372;
  assign T_1350_25 = T_3590;
  assign T_1355_0 = T_3516;
  assign T_1355_1 = T_3616;
  assign T_1355_2 = T_4157;
  assign T_1355_3 = T_4165;
  assign T_1355_4 = T_3916;
  assign T_1355_5 = T_4177;
  assign T_1355_6 = T_4185;
  assign T_1355_7 = T_4193;
  assign T_1355_8 = T_4201;
  assign T_1355_9 = T_3636;
  assign T_1355_10 = T_4213;
  assign T_1355_11 = T_4221;
  assign T_1355_12 = T_3936;
  assign T_1355_13 = T_4235;
  assign T_1355_14 = T_4247;
  assign T_1355_15 = T_4259;
  assign T_1355_16 = T_4273;
  assign T_1355_17 = T_4289;
  assign T_1355_18 = T_4305;
  assign T_1355_19 = T_4321;
  assign T_1355_20 = T_4333;
  assign T_1355_21 = T_4341;
  assign T_1355_22 = T_4351;
  assign T_1355_23 = T_4363;
  assign T_1355_24 = T_4375;
  assign T_1355_25 = T_3596;
  assign T_1360_0 = 1'h1;
  assign T_1360_1 = 1'h1;
  assign T_1360_2 = 1'h1;
  assign T_1360_3 = 1'h1;
  assign T_1360_4 = 1'h1;
  assign T_1360_5 = 1'h1;
  assign T_1360_6 = 1'h1;
  assign T_1360_7 = 1'h1;
  assign T_1360_8 = 1'h1;
  assign T_1360_9 = 1'h1;
  assign T_1360_10 = 1'h1;
  assign T_1360_11 = 1'h1;
  assign T_1360_12 = 1'h1;
  assign T_1360_13 = 1'h1;
  assign T_1360_14 = 1'h1;
  assign T_1360_15 = 1'h1;
  assign T_1360_16 = 1'h1;
  assign T_1360_17 = 1'h1;
  assign T_1360_18 = 1'h1;
  assign T_1360_19 = 1'h1;
  assign T_1360_20 = 1'h1;
  assign T_1360_21 = 1'h1;
  assign T_1360_22 = 1'h1;
  assign T_1360_23 = 1'h1;
  assign T_1360_24 = 1'h1;
  assign T_1360_25 = 1'h1;
  assign T_1365_0 = 1'h1;
  assign T_1365_1 = 1'h1;
  assign T_1365_2 = 1'h1;
  assign T_1365_3 = 1'h1;
  assign T_1365_4 = 1'h1;
  assign T_1365_5 = 1'h1;
  assign T_1365_6 = 1'h1;
  assign T_1365_7 = 1'h1;
  assign T_1365_8 = 1'h1;
  assign T_1365_9 = 1'h1;
  assign T_1365_10 = 1'h1;
  assign T_1365_11 = 1'h1;
  assign T_1365_12 = 1'h1;
  assign T_1365_13 = 1'h1;
  assign T_1365_14 = 1'h1;
  assign T_1365_15 = 1'h1;
  assign T_1365_16 = 1'h1;
  assign T_1365_17 = 1'h1;
  assign T_1365_18 = 1'h1;
  assign T_1365_19 = 1'h1;
  assign T_1365_20 = 1'h1;
  assign T_1365_21 = 1'h1;
  assign T_1365_22 = 1'h1;
  assign T_1365_23 = 1'h1;
  assign T_1365_24 = 1'h1;
  assign T_1365_25 = 1'h1;
  assign T_1370_0 = 1'h1;
  assign T_1370_1 = 1'h1;
  assign T_1370_2 = 1'h1;
  assign T_1370_3 = 1'h1;
  assign T_1370_4 = 1'h1;
  assign T_1370_5 = 1'h1;
  assign T_1370_6 = 1'h1;
  assign T_1370_7 = 1'h1;
  assign T_1370_8 = 1'h1;
  assign T_1370_9 = 1'h1;
  assign T_1370_10 = 1'h1;
  assign T_1370_11 = 1'h1;
  assign T_1370_12 = 1'h1;
  assign T_1370_13 = 1'h1;
  assign T_1370_14 = 1'h1;
  assign T_1370_15 = 1'h1;
  assign T_1370_16 = 1'h1;
  assign T_1370_17 = 1'h1;
  assign T_1370_18 = 1'h1;
  assign T_1370_19 = 1'h1;
  assign T_1370_20 = 1'h1;
  assign T_1370_21 = 1'h1;
  assign T_1370_22 = 1'h1;
  assign T_1370_23 = 1'h1;
  assign T_1370_24 = 1'h1;
  assign T_1370_25 = 1'h1;
  assign T_1375_0 = 1'h1;
  assign T_1375_1 = 1'h1;
  assign T_1375_2 = 1'h1;
  assign T_1375_3 = 1'h1;
  assign T_1375_4 = 1'h1;
  assign T_1375_5 = 1'h1;
  assign T_1375_6 = 1'h1;
  assign T_1375_7 = 1'h1;
  assign T_1375_8 = 1'h1;
  assign T_1375_9 = 1'h1;
  assign T_1375_10 = 1'h1;
  assign T_1375_11 = 1'h1;
  assign T_1375_12 = 1'h1;
  assign T_1375_13 = 1'h1;
  assign T_1375_14 = 1'h1;
  assign T_1375_15 = 1'h1;
  assign T_1375_16 = 1'h1;
  assign T_1375_17 = 1'h1;
  assign T_1375_18 = 1'h1;
  assign T_1375_19 = 1'h1;
  assign T_1375_20 = 1'h1;
  assign T_1375_21 = 1'h1;
  assign T_1375_22 = 1'h1;
  assign T_1375_23 = 1'h1;
  assign T_1375_24 = 1'h1;
  assign T_1375_25 = 1'h1;
  assign T_1380_0 = T_3520;
  assign T_1380_1 = T_3620;
  assign T_1380_2 = T_4159;
  assign T_1380_3 = T_4167;
  assign T_1380_4 = T_3920;
  assign T_1380_5 = T_4179;
  assign T_1380_6 = T_4187;
  assign T_1380_7 = T_4195;
  assign T_1380_8 = T_4203;
  assign T_1380_9 = T_3640;
  assign T_1380_10 = T_4215;
  assign T_1380_11 = T_4223;
  assign T_1380_12 = T_3940;
  assign T_1380_13 = T_4238;
  assign T_1380_14 = T_4250;
  assign T_1380_15 = T_4262;
  assign T_1380_16 = T_4277;
  assign T_1380_17 = T_4293;
  assign T_1380_18 = T_4309;
  assign T_1380_19 = T_4325;
  assign T_1380_20 = T_4335;
  assign T_1380_21 = T_4343;
  assign T_1380_22 = T_4354;
  assign T_1380_23 = T_4366;
  assign T_1380_24 = T_4378;
  assign T_1380_25 = T_3600;
  assign T_1385_0 = T_3526;
  assign T_1385_1 = T_3626;
  assign T_1385_2 = T_4161;
  assign T_1385_3 = T_4169;
  assign T_1385_4 = T_3926;
  assign T_1385_5 = T_4181;
  assign T_1385_6 = T_4189;
  assign T_1385_7 = T_4197;
  assign T_1385_8 = T_4205;
  assign T_1385_9 = T_3646;
  assign T_1385_10 = T_4217;
  assign T_1385_11 = T_4225;
  assign T_1385_12 = T_3946;
  assign T_1385_13 = T_4241;
  assign T_1385_14 = T_4253;
  assign T_1385_15 = T_4265;
  assign T_1385_16 = T_4281;
  assign T_1385_17 = T_4297;
  assign T_1385_18 = T_4313;
  assign T_1385_19 = T_4329;
  assign T_1385_20 = T_4337;
  assign T_1385_21 = T_4345;
  assign T_1385_22 = T_4357;
  assign T_1385_23 = T_4369;
  assign T_1385_24 = T_4381;
  assign T_1385_25 = T_3606;
  assign T_1547 = T_1138_bits_mask[0];
  assign T_1548 = T_1138_bits_mask[1];
  assign T_1549 = T_1138_bits_mask[2];
  assign T_1550 = T_1138_bits_mask[3];
  assign T_1554 = T_1547 ? 8'hff : 8'h0;
  assign T_1558 = T_1548 ? 8'hff : 8'h0;
  assign T_1562 = T_1549 ? 8'hff : 8'h0;
  assign T_1566 = T_1550 ? 8'hff : 8'h0;
  assign T_1567 = {T_1558,T_1554};
  assign T_1568 = {T_1566,T_1562};
  assign T_1569 = {T_1568,T_1567};
  assign T_1593 = T_1569[11:0];
  assign T_1597 = ~ T_1593;
  assign T_1599 = T_1597 == 12'h0;
  assign T_1612 = T_1385_0 & T_1599;
  assign T_1613 = T_1138_bits_data[11:0];
  assign GEN_6 = T_1612 ? T_1613 : ctrl_sck_div;
  assign T_1633 = T_1569[0];
  assign T_1637 = ~ T_1633;
  assign T_1639 = T_1637 == 1'h0;
  assign T_1652 = T_1385_1 & T_1639;
  assign T_1653 = T_1138_bits_data[0];
  assign GEN_7 = T_1652 ? T_1653 : ctrl_cs_dflt_0;
  assign T_1673 = T_1569[7:0];
  assign T_1675 = T_1673 != 8'h0;
  assign T_1677 = ~ T_1673;
  assign T_1679 = T_1677 == 8'h0;
  assign T_1692 = T_1385_2 & T_1679;
  assign T_1693 = T_1138_bits_data[7:0];
  assign GEN_8 = T_1692 ? T_1693 : ctrl_dla_cssck;
  assign T_1713 = T_1569[23:16];
  assign T_1717 = ~ T_1713;
  assign T_1719 = T_1717 == 8'h0;
  assign T_1732 = T_1385_3 & T_1719;
  assign T_1733 = T_1138_bits_data[23:16];
  assign GEN_9 = T_1732 ? T_1733 : ctrl_dla_sckcs;
  assign GEN_210 = {{16'd0}, ctrl_dla_sckcs};
  assign T_1748 = GEN_210 << 16;
  assign GEN_211 = {{16'd0}, ctrl_dla_cssck};
  assign T_1752 = GEN_211 | T_1748;
  assign T_1753 = T_1569[3:0];
  assign T_1757 = ~ T_1753;
  assign T_1759 = T_1757 == 4'h0;
  assign T_1772 = T_1385_4 & T_1759;
  assign T_1773 = T_1138_bits_data[3:0];
  assign GEN_10 = T_1772 ? T_1773 : ctrl_wm_tx;
  assign T_1828 = fifo_io_ip_txwm;
  assign T_1833 = T_1569[1];
  assign T_1837 = ~ T_1833;
  assign T_1839 = T_1837 == 1'h0;
  assign T_1853 = T_1138_bits_data[1];
  assign GEN_212 = {{1'd0}, fifo_io_ip_rxwm};
  assign T_1868 = GEN_212 << 1;
  assign GEN_213 = {{1'd0}, T_1828};
  assign T_1872 = GEN_213 | T_1868;
  assign T_1892 = T_1385_7 & T_1639;
  assign GEN_11 = T_1892 ? T_1653 : ctrl_sck_pha;
  assign T_1932 = T_1385_8 & T_1839;
  assign GEN_12 = T_1932 ? T_1853 : ctrl_sck_pol;
  assign GEN_214 = {{1'd0}, ctrl_sck_pol};
  assign T_1948 = GEN_214 << 1;
  assign GEN_215 = {{1'd0}, ctrl_sck_pha};
  assign T_1952 = GEN_215 | T_1948;
  assign T_1953 = T_1569[1:0];
  assign T_1957 = ~ T_1953;
  assign T_1959 = T_1957 == 2'h0;
  assign T_1972 = T_1385_9 & T_1959;
  assign T_1973 = T_1138_bits_data[1:0];
  assign GEN_13 = T_1972 ? T_1973 : ctrl_cs_mode;
  assign T_2012 = T_1385_10 & T_1639;
  assign GEN_14 = T_2012 ? T_1653 : ie_txwm;
  assign T_2052 = T_1385_11 & T_1839;
  assign GEN_15 = T_2052 ? T_1853 : ie_rxwm;
  assign GEN_216 = {{1'd0}, ie_rxwm};
  assign T_2068 = GEN_216 << 1;
  assign GEN_217 = {{1'd0}, ie_txwm};
  assign T_2072 = GEN_217 | T_2068;
  assign T_2092 = T_1385_12 & T_1759;
  assign GEN_16 = T_2092 ? T_1773 : ctrl_wm_rx;
  assign T_2132 = T_1385_13 & T_1679;
  assign GEN_218 = {{31'd0}, T_1036};
  assign T_2228 = GEN_218 << 31;
  assign T_2252 = T_1385_16 & T_1959;
  assign GEN_17 = T_2252 ? T_1973 : ctrl_fmt_proto;
  assign T_2273 = T_1569[2];
  assign T_2277 = ~ T_2273;
  assign T_2279 = T_2277 == 1'h0;
  assign T_2292 = T_1385_17 & T_2279;
  assign T_2293 = T_1138_bits_data[2];
  assign GEN_18 = T_2292 ? T_2293 : ctrl_fmt_endian;
  assign GEN_219 = {{2'd0}, ctrl_fmt_endian};
  assign T_2308 = GEN_219 << 2;
  assign GEN_220 = {{1'd0}, ctrl_fmt_proto};
  assign T_2312 = GEN_220 | T_2308;
  assign T_2313 = T_1569[3];
  assign T_2317 = ~ T_2313;
  assign T_2319 = T_2317 == 1'h0;
  assign T_2332 = T_1385_18 & T_2319;
  assign T_2333 = T_1138_bits_data[3];
  assign GEN_19 = T_2332 ? T_2333 : ctrl_fmt_iodir;
  assign GEN_221 = {{3'd0}, ctrl_fmt_iodir};
  assign T_2348 = GEN_221 << 3;
  assign GEN_222 = {{1'd0}, T_2312};
  assign T_2352 = GEN_222 | T_2348;
  assign T_2353 = T_1569[19:16];
  assign T_2357 = ~ T_2353;
  assign T_2359 = T_2357 == 4'h0;
  assign T_2372 = T_1385_19 & T_2359;
  assign T_2373 = T_1138_bits_data[19:16];
  assign GEN_20 = T_2372 ? T_2373 : ctrl_fmt_len;
  assign GEN_223 = {{16'd0}, ctrl_fmt_len};
  assign T_2388 = GEN_223 << 16;
  assign GEN_224 = {{16'd0}, T_2352};
  assign T_2392 = GEN_224 | T_2388;
  assign T_2412 = T_1385_20 & T_1679;
  assign GEN_21 = T_2412 ? T_1693 : ctrl_dla_intercs;
  assign T_2452 = T_1385_21 & T_1719;
  assign GEN_22 = T_2452 ? T_1733 : ctrl_dla_interxfr;
  assign GEN_225 = {{16'd0}, ctrl_dla_interxfr};
  assign T_2468 = GEN_225 << 16;
  assign GEN_226 = {{16'd0}, ctrl_dla_intercs};
  assign T_2472 = GEN_226 | T_2468;
  assign T_2488 = T_1380_22 & T_1675;
  assign T_2508 = fifo_io_rx_bits;
  assign T_2552 = {{23'd0}, T_2508};
  assign GEN_227 = {{31'd0}, T_1039};
  assign T_2588 = GEN_227 << 31;
  assign GEN_228 = {{1'd0}, T_2552};
  assign T_2592 = GEN_228 | T_2588;
  assign T_2612 = T_1385_25 & T_1639;
  assign GEN_23 = T_2612 ? T_1653 : ctrl_cs_id;
  assign T_2634 = T_1225 == 1'h0;
  assign T_2636 = T_2634 | T_1360_0;
  assign T_2638 = T_1270 == 1'h0;
  assign T_2639 = T_1360_8 & T_1360_7;
  assign T_2641 = T_2638 | T_2639;
  assign T_2649 = T_1342 == 1'h0;
  assign T_2651 = T_2649 | T_1360_25;
  assign T_2653 = T_1234 == 1'h0;
  assign T_2655 = T_2653 | T_1360_1;
  assign T_2657 = T_1279 == 1'h0;
  assign T_2659 = T_2657 | T_1360_9;
  assign T_2670 = T_1243 == 1'h0;
  assign T_2671 = T_1360_3 & T_1360_2;
  assign T_2673 = T_2670 | T_2671;
  assign T_2675 = T_1324 == 1'h0;
  assign T_2676 = T_1360_21 & T_1360_20;
  assign T_2678 = T_2675 | T_2676;
  assign T_2692 = T_1315 == 1'h0;
  assign T_2693 = T_1360_19 & T_1360_18;
  assign T_2694 = T_2693 & T_1360_17;
  assign T_2695 = T_2694 & T_1360_16;
  assign T_2697 = T_2692 | T_2695;
  assign T_2702 = T_1306 == 1'h0;
  assign T_2703 = T_1360_15 & T_1360_14;
  assign T_2704 = T_2703 & T_1360_13;
  assign T_2706 = T_2702 | T_2704;
  assign T_2708 = T_1333 == 1'h0;
  assign T_2709 = T_1360_24 & T_1360_23;
  assign T_2710 = T_2709 & T_1360_22;
  assign T_2712 = T_2708 | T_2710;
  assign T_2714 = T_1252 == 1'h0;
  assign T_2716 = T_2714 | T_1360_4;
  assign T_2718 = T_1297 == 1'h0;
  assign T_2720 = T_2718 | T_1360_12;
  assign T_2740 = T_1288 == 1'h0;
  assign T_2741 = T_1360_11 & T_1360_10;
  assign T_2743 = T_2740 | T_2741;
  assign T_2745 = T_1261 == 1'h0;
  assign T_2746 = T_1360_6 & T_1360_5;
  assign T_2748 = T_2745 | T_2746;
  assign T_2790_0 = T_2636;
  assign T_2790_1 = T_2641;
  assign T_2790_2 = 1'h1;
  assign T_2790_3 = 1'h1;
  assign T_2790_4 = T_2651;
  assign T_2790_5 = T_2655;
  assign T_2790_6 = T_2659;
  assign T_2790_7 = 1'h1;
  assign T_2790_8 = 1'h1;
  assign T_2790_9 = 1'h1;
  assign T_2790_10 = T_2673;
  assign T_2790_11 = T_2678;
  assign T_2790_12 = 1'h1;
  assign T_2790_13 = 1'h1;
  assign T_2790_14 = 1'h1;
  assign T_2790_15 = 1'h1;
  assign T_2790_16 = T_2697;
  assign T_2790_17 = 1'h1;
  assign T_2790_18 = T_2706;
  assign T_2790_19 = T_2712;
  assign T_2790_20 = T_2716;
  assign T_2790_21 = T_2720;
  assign T_2790_22 = 1'h1;
  assign T_2790_23 = 1'h1;
  assign T_2790_24 = 1'h1;
  assign T_2790_25 = 1'h1;
  assign T_2790_26 = 1'h1;
  assign T_2790_27 = 1'h1;
  assign T_2790_28 = T_2743;
  assign T_2790_29 = T_2748;
  assign T_2790_30 = 1'h1;
  assign T_2790_31 = 1'h1;
  assign T_2828 = T_2634 | T_1365_0;
  assign T_2831 = T_1365_8 & T_1365_7;
  assign T_2833 = T_2638 | T_2831;
  assign T_2843 = T_2649 | T_1365_25;
  assign T_2847 = T_2653 | T_1365_1;
  assign T_2851 = T_2657 | T_1365_9;
  assign T_2863 = T_1365_3 & T_1365_2;
  assign T_2865 = T_2670 | T_2863;
  assign T_2868 = T_1365_21 & T_1365_20;
  assign T_2870 = T_2675 | T_2868;
  assign T_2885 = T_1365_19 & T_1365_18;
  assign T_2886 = T_2885 & T_1365_17;
  assign T_2887 = T_2886 & T_1365_16;
  assign T_2889 = T_2692 | T_2887;
  assign T_2895 = T_1365_15 & T_1365_14;
  assign T_2896 = T_2895 & T_1365_13;
  assign T_2898 = T_2702 | T_2896;
  assign T_2901 = T_1365_24 & T_1365_23;
  assign T_2902 = T_2901 & T_1365_22;
  assign T_2904 = T_2708 | T_2902;
  assign T_2908 = T_2714 | T_1365_4;
  assign T_2912 = T_2718 | T_1365_12;
  assign T_2933 = T_1365_11 & T_1365_10;
  assign T_2935 = T_2740 | T_2933;
  assign T_2938 = T_1365_6 & T_1365_5;
  assign T_2940 = T_2745 | T_2938;
  assign T_2982_0 = T_2828;
  assign T_2982_1 = T_2833;
  assign T_2982_2 = 1'h1;
  assign T_2982_3 = 1'h1;
  assign T_2982_4 = T_2843;
  assign T_2982_5 = T_2847;
  assign T_2982_6 = T_2851;
  assign T_2982_7 = 1'h1;
  assign T_2982_8 = 1'h1;
  assign T_2982_9 = 1'h1;
  assign T_2982_10 = T_2865;
  assign T_2982_11 = T_2870;
  assign T_2982_12 = 1'h1;
  assign T_2982_13 = 1'h1;
  assign T_2982_14 = 1'h1;
  assign T_2982_15 = 1'h1;
  assign T_2982_16 = T_2889;
  assign T_2982_17 = 1'h1;
  assign T_2982_18 = T_2898;
  assign T_2982_19 = T_2904;
  assign T_2982_20 = T_2908;
  assign T_2982_21 = T_2912;
  assign T_2982_22 = 1'h1;
  assign T_2982_23 = 1'h1;
  assign T_2982_24 = 1'h1;
  assign T_2982_25 = 1'h1;
  assign T_2982_26 = 1'h1;
  assign T_2982_27 = 1'h1;
  assign T_2982_28 = T_2935;
  assign T_2982_29 = T_2940;
  assign T_2982_30 = 1'h1;
  assign T_2982_31 = 1'h1;
  assign T_3020 = T_2634 | T_1370_0;
  assign T_3023 = T_1370_8 & T_1370_7;
  assign T_3025 = T_2638 | T_3023;
  assign T_3035 = T_2649 | T_1370_25;
  assign T_3039 = T_2653 | T_1370_1;
  assign T_3043 = T_2657 | T_1370_9;
  assign T_3055 = T_1370_3 & T_1370_2;
  assign T_3057 = T_2670 | T_3055;
  assign T_3060 = T_1370_21 & T_1370_20;
  assign T_3062 = T_2675 | T_3060;
  assign T_3077 = T_1370_19 & T_1370_18;
  assign T_3078 = T_3077 & T_1370_17;
  assign T_3079 = T_3078 & T_1370_16;
  assign T_3081 = T_2692 | T_3079;
  assign T_3087 = T_1370_15 & T_1370_14;
  assign T_3088 = T_3087 & T_1370_13;
  assign T_3090 = T_2702 | T_3088;
  assign T_3093 = T_1370_24 & T_1370_23;
  assign T_3094 = T_3093 & T_1370_22;
  assign T_3096 = T_2708 | T_3094;
  assign T_3100 = T_2714 | T_1370_4;
  assign T_3104 = T_2718 | T_1370_12;
  assign T_3125 = T_1370_11 & T_1370_10;
  assign T_3127 = T_2740 | T_3125;
  assign T_3130 = T_1370_6 & T_1370_5;
  assign T_3132 = T_2745 | T_3130;
  assign T_3174_0 = T_3020;
  assign T_3174_1 = T_3025;
  assign T_3174_2 = 1'h1;
  assign T_3174_3 = 1'h1;
  assign T_3174_4 = T_3035;
  assign T_3174_5 = T_3039;
  assign T_3174_6 = T_3043;
  assign T_3174_7 = 1'h1;
  assign T_3174_8 = 1'h1;
  assign T_3174_9 = 1'h1;
  assign T_3174_10 = T_3057;
  assign T_3174_11 = T_3062;
  assign T_3174_12 = 1'h1;
  assign T_3174_13 = 1'h1;
  assign T_3174_14 = 1'h1;
  assign T_3174_15 = 1'h1;
  assign T_3174_16 = T_3081;
  assign T_3174_17 = 1'h1;
  assign T_3174_18 = T_3090;
  assign T_3174_19 = T_3096;
  assign T_3174_20 = T_3100;
  assign T_3174_21 = T_3104;
  assign T_3174_22 = 1'h1;
  assign T_3174_23 = 1'h1;
  assign T_3174_24 = 1'h1;
  assign T_3174_25 = 1'h1;
  assign T_3174_26 = 1'h1;
  assign T_3174_27 = 1'h1;
  assign T_3174_28 = T_3127;
  assign T_3174_29 = T_3132;
  assign T_3174_30 = 1'h1;
  assign T_3174_31 = 1'h1;
  assign T_3212 = T_2634 | T_1375_0;
  assign T_3215 = T_1375_8 & T_1375_7;
  assign T_3217 = T_2638 | T_3215;
  assign T_3227 = T_2649 | T_1375_25;
  assign T_3231 = T_2653 | T_1375_1;
  assign T_3235 = T_2657 | T_1375_9;
  assign T_3247 = T_1375_3 & T_1375_2;
  assign T_3249 = T_2670 | T_3247;
  assign T_3252 = T_1375_21 & T_1375_20;
  assign T_3254 = T_2675 | T_3252;
  assign T_3269 = T_1375_19 & T_1375_18;
  assign T_3270 = T_3269 & T_1375_17;
  assign T_3271 = T_3270 & T_1375_16;
  assign T_3273 = T_2692 | T_3271;
  assign T_3279 = T_1375_15 & T_1375_14;
  assign T_3280 = T_3279 & T_1375_13;
  assign T_3282 = T_2702 | T_3280;
  assign T_3285 = T_1375_24 & T_1375_23;
  assign T_3286 = T_3285 & T_1375_22;
  assign T_3288 = T_2708 | T_3286;
  assign T_3292 = T_2714 | T_1375_4;
  assign T_3296 = T_2718 | T_1375_12;
  assign T_3317 = T_1375_11 & T_1375_10;
  assign T_3319 = T_2740 | T_3317;
  assign T_3322 = T_1375_6 & T_1375_5;
  assign T_3324 = T_2745 | T_3322;
  assign T_3366_0 = T_3212;
  assign T_3366_1 = T_3217;
  assign T_3366_2 = 1'h1;
  assign T_3366_3 = 1'h1;
  assign T_3366_4 = T_3227;
  assign T_3366_5 = T_3231;
  assign T_3366_6 = T_3235;
  assign T_3366_7 = 1'h1;
  assign T_3366_8 = 1'h1;
  assign T_3366_9 = 1'h1;
  assign T_3366_10 = T_3249;
  assign T_3366_11 = T_3254;
  assign T_3366_12 = 1'h1;
  assign T_3366_13 = 1'h1;
  assign T_3366_14 = 1'h1;
  assign T_3366_15 = 1'h1;
  assign T_3366_16 = T_3273;
  assign T_3366_17 = 1'h1;
  assign T_3366_18 = T_3282;
  assign T_3366_19 = T_3288;
  assign T_3366_20 = T_3292;
  assign T_3366_21 = T_3296;
  assign T_3366_22 = 1'h1;
  assign T_3366_23 = 1'h1;
  assign T_3366_24 = 1'h1;
  assign T_3366_25 = 1'h1;
  assign T_3366_26 = 1'h1;
  assign T_3366_27 = 1'h1;
  assign T_3366_28 = T_3319;
  assign T_3366_29 = T_3324;
  assign T_3366_30 = 1'h1;
  assign T_3366_31 = 1'h1;
  assign T_3401 = T_1138_bits_index[0];
  assign T_3402 = T_1138_bits_index[1];
  assign T_3403 = T_1138_bits_index[2];
  assign T_3404 = T_1138_bits_index[3];
  assign T_3405 = T_1138_bits_index[4];
  assign T_3411 = {T_3402,T_3401};
  assign T_3412 = {T_3405,T_3404};
  assign T_3413 = {T_3412,T_3403};
  assign T_3414 = {T_3413,T_3411};
  assign GEN_0 = GEN_54;
  assign GEN_24 = 5'h1 == T_3414 ? T_2790_1 : T_2790_0;
  assign GEN_25 = 5'h2 == T_3414 ? T_2790_2 : GEN_24;
  assign GEN_26 = 5'h3 == T_3414 ? T_2790_3 : GEN_25;
  assign GEN_27 = 5'h4 == T_3414 ? T_2790_4 : GEN_26;
  assign GEN_28 = 5'h5 == T_3414 ? T_2790_5 : GEN_27;
  assign GEN_29 = 5'h6 == T_3414 ? T_2790_6 : GEN_28;
  assign GEN_30 = 5'h7 == T_3414 ? T_2790_7 : GEN_29;
  assign GEN_31 = 5'h8 == T_3414 ? T_2790_8 : GEN_30;
  assign GEN_32 = 5'h9 == T_3414 ? T_2790_9 : GEN_31;
  assign GEN_33 = 5'ha == T_3414 ? T_2790_10 : GEN_32;
  assign GEN_34 = 5'hb == T_3414 ? T_2790_11 : GEN_33;
  assign GEN_35 = 5'hc == T_3414 ? T_2790_12 : GEN_34;
  assign GEN_36 = 5'hd == T_3414 ? T_2790_13 : GEN_35;
  assign GEN_37 = 5'he == T_3414 ? T_2790_14 : GEN_36;
  assign GEN_38 = 5'hf == T_3414 ? T_2790_15 : GEN_37;
  assign GEN_39 = 5'h10 == T_3414 ? T_2790_16 : GEN_38;
  assign GEN_40 = 5'h11 == T_3414 ? T_2790_17 : GEN_39;
  assign GEN_41 = 5'h12 == T_3414 ? T_2790_18 : GEN_40;
  assign GEN_42 = 5'h13 == T_3414 ? T_2790_19 : GEN_41;
  assign GEN_43 = 5'h14 == T_3414 ? T_2790_20 : GEN_42;
  assign GEN_44 = 5'h15 == T_3414 ? T_2790_21 : GEN_43;
  assign GEN_45 = 5'h16 == T_3414 ? T_2790_22 : GEN_44;
  assign GEN_46 = 5'h17 == T_3414 ? T_2790_23 : GEN_45;
  assign GEN_47 = 5'h18 == T_3414 ? T_2790_24 : GEN_46;
  assign GEN_48 = 5'h19 == T_3414 ? T_2790_25 : GEN_47;
  assign GEN_49 = 5'h1a == T_3414 ? T_2790_26 : GEN_48;
  assign GEN_50 = 5'h1b == T_3414 ? T_2790_27 : GEN_49;
  assign GEN_51 = 5'h1c == T_3414 ? T_2790_28 : GEN_50;
  assign GEN_52 = 5'h1d == T_3414 ? T_2790_29 : GEN_51;
  assign GEN_53 = 5'h1e == T_3414 ? T_2790_30 : GEN_52;
  assign GEN_54 = 5'h1f == T_3414 ? T_2790_31 : GEN_53;
  assign GEN_1 = GEN_85;
  assign GEN_55 = 5'h1 == T_3414 ? T_2982_1 : T_2982_0;
  assign GEN_56 = 5'h2 == T_3414 ? T_2982_2 : GEN_55;
  assign GEN_57 = 5'h3 == T_3414 ? T_2982_3 : GEN_56;
  assign GEN_58 = 5'h4 == T_3414 ? T_2982_4 : GEN_57;
  assign GEN_59 = 5'h5 == T_3414 ? T_2982_5 : GEN_58;
  assign GEN_60 = 5'h6 == T_3414 ? T_2982_6 : GEN_59;
  assign GEN_61 = 5'h7 == T_3414 ? T_2982_7 : GEN_60;
  assign GEN_62 = 5'h8 == T_3414 ? T_2982_8 : GEN_61;
  assign GEN_63 = 5'h9 == T_3414 ? T_2982_9 : GEN_62;
  assign GEN_64 = 5'ha == T_3414 ? T_2982_10 : GEN_63;
  assign GEN_65 = 5'hb == T_3414 ? T_2982_11 : GEN_64;
  assign GEN_66 = 5'hc == T_3414 ? T_2982_12 : GEN_65;
  assign GEN_67 = 5'hd == T_3414 ? T_2982_13 : GEN_66;
  assign GEN_68 = 5'he == T_3414 ? T_2982_14 : GEN_67;
  assign GEN_69 = 5'hf == T_3414 ? T_2982_15 : GEN_68;
  assign GEN_70 = 5'h10 == T_3414 ? T_2982_16 : GEN_69;
  assign GEN_71 = 5'h11 == T_3414 ? T_2982_17 : GEN_70;
  assign GEN_72 = 5'h12 == T_3414 ? T_2982_18 : GEN_71;
  assign GEN_73 = 5'h13 == T_3414 ? T_2982_19 : GEN_72;
  assign GEN_74 = 5'h14 == T_3414 ? T_2982_20 : GEN_73;
  assign GEN_75 = 5'h15 == T_3414 ? T_2982_21 : GEN_74;
  assign GEN_76 = 5'h16 == T_3414 ? T_2982_22 : GEN_75;
  assign GEN_77 = 5'h17 == T_3414 ? T_2982_23 : GEN_76;
  assign GEN_78 = 5'h18 == T_3414 ? T_2982_24 : GEN_77;
  assign GEN_79 = 5'h19 == T_3414 ? T_2982_25 : GEN_78;
  assign GEN_80 = 5'h1a == T_3414 ? T_2982_26 : GEN_79;
  assign GEN_81 = 5'h1b == T_3414 ? T_2982_27 : GEN_80;
  assign GEN_82 = 5'h1c == T_3414 ? T_2982_28 : GEN_81;
  assign GEN_83 = 5'h1d == T_3414 ? T_2982_29 : GEN_82;
  assign GEN_84 = 5'h1e == T_3414 ? T_2982_30 : GEN_83;
  assign GEN_85 = 5'h1f == T_3414 ? T_2982_31 : GEN_84;
  assign T_3431 = T_1138_bits_read ? GEN_0 : GEN_1;
  assign GEN_2 = GEN_116;
  assign GEN_86 = 5'h1 == T_3414 ? T_3174_1 : T_3174_0;
  assign GEN_87 = 5'h2 == T_3414 ? T_3174_2 : GEN_86;
  assign GEN_88 = 5'h3 == T_3414 ? T_3174_3 : GEN_87;
  assign GEN_89 = 5'h4 == T_3414 ? T_3174_4 : GEN_88;
  assign GEN_90 = 5'h5 == T_3414 ? T_3174_5 : GEN_89;
  assign GEN_91 = 5'h6 == T_3414 ? T_3174_6 : GEN_90;
  assign GEN_92 = 5'h7 == T_3414 ? T_3174_7 : GEN_91;
  assign GEN_93 = 5'h8 == T_3414 ? T_3174_8 : GEN_92;
  assign GEN_94 = 5'h9 == T_3414 ? T_3174_9 : GEN_93;
  assign GEN_95 = 5'ha == T_3414 ? T_3174_10 : GEN_94;
  assign GEN_96 = 5'hb == T_3414 ? T_3174_11 : GEN_95;
  assign GEN_97 = 5'hc == T_3414 ? T_3174_12 : GEN_96;
  assign GEN_98 = 5'hd == T_3414 ? T_3174_13 : GEN_97;
  assign GEN_99 = 5'he == T_3414 ? T_3174_14 : GEN_98;
  assign GEN_100 = 5'hf == T_3414 ? T_3174_15 : GEN_99;
  assign GEN_101 = 5'h10 == T_3414 ? T_3174_16 : GEN_100;
  assign GEN_102 = 5'h11 == T_3414 ? T_3174_17 : GEN_101;
  assign GEN_103 = 5'h12 == T_3414 ? T_3174_18 : GEN_102;
  assign GEN_104 = 5'h13 == T_3414 ? T_3174_19 : GEN_103;
  assign GEN_105 = 5'h14 == T_3414 ? T_3174_20 : GEN_104;
  assign GEN_106 = 5'h15 == T_3414 ? T_3174_21 : GEN_105;
  assign GEN_107 = 5'h16 == T_3414 ? T_3174_22 : GEN_106;
  assign GEN_108 = 5'h17 == T_3414 ? T_3174_23 : GEN_107;
  assign GEN_109 = 5'h18 == T_3414 ? T_3174_24 : GEN_108;
  assign GEN_110 = 5'h19 == T_3414 ? T_3174_25 : GEN_109;
  assign GEN_111 = 5'h1a == T_3414 ? T_3174_26 : GEN_110;
  assign GEN_112 = 5'h1b == T_3414 ? T_3174_27 : GEN_111;
  assign GEN_113 = 5'h1c == T_3414 ? T_3174_28 : GEN_112;
  assign GEN_114 = 5'h1d == T_3414 ? T_3174_29 : GEN_113;
  assign GEN_115 = 5'h1e == T_3414 ? T_3174_30 : GEN_114;
  assign GEN_116 = 5'h1f == T_3414 ? T_3174_31 : GEN_115;
  assign GEN_3 = GEN_147;
  assign GEN_117 = 5'h1 == T_3414 ? T_3366_1 : T_3366_0;
  assign GEN_118 = 5'h2 == T_3414 ? T_3366_2 : GEN_117;
  assign GEN_119 = 5'h3 == T_3414 ? T_3366_3 : GEN_118;
  assign GEN_120 = 5'h4 == T_3414 ? T_3366_4 : GEN_119;
  assign GEN_121 = 5'h5 == T_3414 ? T_3366_5 : GEN_120;
  assign GEN_122 = 5'h6 == T_3414 ? T_3366_6 : GEN_121;
  assign GEN_123 = 5'h7 == T_3414 ? T_3366_7 : GEN_122;
  assign GEN_124 = 5'h8 == T_3414 ? T_3366_8 : GEN_123;
  assign GEN_125 = 5'h9 == T_3414 ? T_3366_9 : GEN_124;
  assign GEN_126 = 5'ha == T_3414 ? T_3366_10 : GEN_125;
  assign GEN_127 = 5'hb == T_3414 ? T_3366_11 : GEN_126;
  assign GEN_128 = 5'hc == T_3414 ? T_3366_12 : GEN_127;
  assign GEN_129 = 5'hd == T_3414 ? T_3366_13 : GEN_128;
  assign GEN_130 = 5'he == T_3414 ? T_3366_14 : GEN_129;
  assign GEN_131 = 5'hf == T_3414 ? T_3366_15 : GEN_130;
  assign GEN_132 = 5'h10 == T_3414 ? T_3366_16 : GEN_131;
  assign GEN_133 = 5'h11 == T_3414 ? T_3366_17 : GEN_132;
  assign GEN_134 = 5'h12 == T_3414 ? T_3366_18 : GEN_133;
  assign GEN_135 = 5'h13 == T_3414 ? T_3366_19 : GEN_134;
  assign GEN_136 = 5'h14 == T_3414 ? T_3366_20 : GEN_135;
  assign GEN_137 = 5'h15 == T_3414 ? T_3366_21 : GEN_136;
  assign GEN_138 = 5'h16 == T_3414 ? T_3366_22 : GEN_137;
  assign GEN_139 = 5'h17 == T_3414 ? T_3366_23 : GEN_138;
  assign GEN_140 = 5'h18 == T_3414 ? T_3366_24 : GEN_139;
  assign GEN_141 = 5'h19 == T_3414 ? T_3366_25 : GEN_140;
  assign GEN_142 = 5'h1a == T_3414 ? T_3366_26 : GEN_141;
  assign GEN_143 = 5'h1b == T_3414 ? T_3366_27 : GEN_142;
  assign GEN_144 = 5'h1c == T_3414 ? T_3366_28 : GEN_143;
  assign GEN_145 = 5'h1d == T_3414 ? T_3366_29 : GEN_144;
  assign GEN_146 = 5'h1e == T_3414 ? T_3366_30 : GEN_145;
  assign GEN_147 = 5'h1f == T_3414 ? T_3366_31 : GEN_146;
  assign T_3434 = T_1138_bits_read ? GEN_2 : GEN_3;
  assign T_3435 = T_1138_ready & T_3431;
  assign T_3436 = T_1063_valid & T_3431;
  assign T_3437 = T_1102_ready & T_3434;
  assign T_3438 = T_1138_valid & T_3434;
  assign T_3440 = 32'h1 << T_3414;
  assign T_3441 = {T_1270,T_1225};
  assign T_3443 = {2'h3,T_3441};
  assign T_3444 = {T_1234,T_1342};
  assign T_3445 = {1'h1,T_1279};
  assign T_3446 = {T_3445,T_3444};
  assign T_3447 = {T_3446,T_3443};
  assign T_3449 = {T_1324,T_1243};
  assign T_3450 = {T_3449,2'h3};
  assign T_3454 = {4'hf,T_3450};
  assign T_3455 = {T_3454,T_3447};
  assign T_3456 = {1'h1,T_1315};
  assign T_3457 = {T_1333,T_1306};
  assign T_3458 = {T_3457,T_3456};
  assign T_3459 = {T_1297,T_1252};
  assign T_3461 = {2'h3,T_3459};
  assign T_3462 = {T_3461,T_3458};
  assign T_3466 = {T_1261,T_1288};
  assign T_3468 = {2'h3,T_3466};
  assign T_3469 = {T_3468,4'hf};
  assign T_3470 = {T_3469,T_3462};
  assign T_3471 = {T_3470,T_3455};
  assign T_3472 = T_3440 & T_3471;
  assign T_3507 = T_1063_valid & T_1138_ready;
  assign T_3508 = T_3507 & T_1138_bits_read;
  assign T_3509 = T_3472[0];
  assign T_3510 = T_3508 & T_3509;
  assign T_3513 = T_1138_bits_read == 1'h0;
  assign T_3514 = T_3507 & T_3513;
  assign T_3516 = T_3514 & T_3509;
  assign T_3517 = T_1138_valid & T_1102_ready;
  assign T_3518 = T_3517 & T_1138_bits_read;
  assign T_3520 = T_3518 & T_3509;
  assign T_3524 = T_3517 & T_3513;
  assign T_3526 = T_3524 & T_3509;
  assign T_3529 = T_3472[1];
  assign T_3530 = T_3508 & T_3529;
  assign T_3536 = T_3514 & T_3529;
  assign T_3540 = T_3518 & T_3529;
  assign T_3546 = T_3524 & T_3529;
  assign T_3589 = T_3472[4];
  assign T_3590 = T_3508 & T_3589;
  assign T_3596 = T_3514 & T_3589;
  assign T_3600 = T_3518 & T_3589;
  assign T_3606 = T_3524 & T_3589;
  assign T_3609 = T_3472[5];
  assign T_3610 = T_3508 & T_3609;
  assign T_3616 = T_3514 & T_3609;
  assign T_3620 = T_3518 & T_3609;
  assign T_3626 = T_3524 & T_3609;
  assign T_3629 = T_3472[6];
  assign T_3630 = T_3508 & T_3629;
  assign T_3636 = T_3514 & T_3629;
  assign T_3640 = T_3518 & T_3629;
  assign T_3646 = T_3524 & T_3629;
  assign T_3709 = T_3472[10];
  assign T_3710 = T_3508 & T_3709;
  assign T_3716 = T_3514 & T_3709;
  assign T_3720 = T_3518 & T_3709;
  assign T_3726 = T_3524 & T_3709;
  assign T_3729 = T_3472[11];
  assign T_3730 = T_3508 & T_3729;
  assign T_3736 = T_3514 & T_3729;
  assign T_3740 = T_3518 & T_3729;
  assign T_3746 = T_3524 & T_3729;
  assign T_3829 = T_3472[16];
  assign T_3830 = T_3508 & T_3829;
  assign T_3836 = T_3514 & T_3829;
  assign T_3840 = T_3518 & T_3829;
  assign T_3846 = T_3524 & T_3829;
  assign T_3869 = T_3472[18];
  assign T_3870 = T_3508 & T_3869;
  assign T_3876 = T_3514 & T_3869;
  assign T_3880 = T_3518 & T_3869;
  assign T_3886 = T_3524 & T_3869;
  assign T_3889 = T_3472[19];
  assign T_3890 = T_3508 & T_3889;
  assign T_3896 = T_3514 & T_3889;
  assign T_3900 = T_3518 & T_3889;
  assign T_3906 = T_3524 & T_3889;
  assign T_3909 = T_3472[20];
  assign T_3910 = T_3508 & T_3909;
  assign T_3916 = T_3514 & T_3909;
  assign T_3920 = T_3518 & T_3909;
  assign T_3926 = T_3524 & T_3909;
  assign T_3929 = T_3472[21];
  assign T_3930 = T_3508 & T_3929;
  assign T_3936 = T_3514 & T_3929;
  assign T_3940 = T_3518 & T_3929;
  assign T_3946 = T_3524 & T_3929;
  assign T_4069 = T_3472[28];
  assign T_4070 = T_3508 & T_4069;
  assign T_4076 = T_3514 & T_4069;
  assign T_4080 = T_3518 & T_4069;
  assign T_4086 = T_3524 & T_4069;
  assign T_4089 = T_3472[29];
  assign T_4090 = T_3508 & T_4089;
  assign T_4096 = T_3514 & T_4089;
  assign T_4100 = T_3518 & T_4089;
  assign T_4106 = T_3524 & T_4089;
  assign T_4155 = T_3710 & T_1360_3;
  assign T_4157 = T_3716 & T_1365_3;
  assign T_4159 = T_3720 & T_1370_3;
  assign T_4161 = T_3726 & T_1375_3;
  assign T_4163 = T_3710 & T_1360_2;
  assign T_4165 = T_3716 & T_1365_2;
  assign T_4167 = T_3720 & T_1370_2;
  assign T_4169 = T_3726 & T_1375_2;
  assign T_4175 = T_4090 & T_1360_6;
  assign T_4177 = T_4096 & T_1365_6;
  assign T_4179 = T_4100 & T_1370_6;
  assign T_4181 = T_4106 & T_1375_6;
  assign T_4183 = T_4090 & T_1360_5;
  assign T_4185 = T_4096 & T_1365_5;
  assign T_4187 = T_4100 & T_1370_5;
  assign T_4189 = T_4106 & T_1375_5;
  assign T_4191 = T_3530 & T_1360_8;
  assign T_4193 = T_3536 & T_1365_8;
  assign T_4195 = T_3540 & T_1370_8;
  assign T_4197 = T_3546 & T_1375_8;
  assign T_4199 = T_3530 & T_1360_7;
  assign T_4201 = T_3536 & T_1365_7;
  assign T_4203 = T_3540 & T_1370_7;
  assign T_4205 = T_3546 & T_1375_7;
  assign T_4211 = T_4070 & T_1360_11;
  assign T_4213 = T_4076 & T_1365_11;
  assign T_4215 = T_4080 & T_1370_11;
  assign T_4217 = T_4086 & T_1375_11;
  assign T_4219 = T_4070 & T_1360_10;
  assign T_4221 = T_4076 & T_1365_10;
  assign T_4223 = T_4080 & T_1370_10;
  assign T_4225 = T_4086 & T_1375_10;
  assign T_4231 = T_3870 & T_1360_15;
  assign T_4232 = T_4231 & T_1360_14;
  assign T_4234 = T_3876 & T_1365_15;
  assign T_4235 = T_4234 & T_1365_14;
  assign T_4237 = T_3880 & T_1370_15;
  assign T_4238 = T_4237 & T_1370_14;
  assign T_4240 = T_3886 & T_1375_15;
  assign T_4241 = T_4240 & T_1375_14;
  assign T_4244 = T_4231 & T_1360_13;
  assign T_4247 = T_4234 & T_1365_13;
  assign T_4250 = T_4237 & T_1370_13;
  assign T_4253 = T_4240 & T_1375_13;
  assign T_4255 = T_3870 & T_1360_14;
  assign T_4256 = T_4255 & T_1360_13;
  assign T_4258 = T_3876 & T_1365_14;
  assign T_4259 = T_4258 & T_1365_13;
  assign T_4261 = T_3880 & T_1370_14;
  assign T_4262 = T_4261 & T_1370_13;
  assign T_4264 = T_3886 & T_1375_14;
  assign T_4265 = T_4264 & T_1375_13;
  assign T_4267 = T_3830 & T_1360_19;
  assign T_4268 = T_4267 & T_1360_18;
  assign T_4269 = T_4268 & T_1360_17;
  assign T_4271 = T_3836 & T_1365_19;
  assign T_4272 = T_4271 & T_1365_18;
  assign T_4273 = T_4272 & T_1365_17;
  assign T_4275 = T_3840 & T_1370_19;
  assign T_4276 = T_4275 & T_1370_18;
  assign T_4277 = T_4276 & T_1370_17;
  assign T_4279 = T_3846 & T_1375_19;
  assign T_4280 = T_4279 & T_1375_18;
  assign T_4281 = T_4280 & T_1375_17;
  assign T_4285 = T_4268 & T_1360_16;
  assign T_4289 = T_4272 & T_1365_16;
  assign T_4293 = T_4276 & T_1370_16;
  assign T_4297 = T_4280 & T_1375_16;
  assign T_4300 = T_4267 & T_1360_17;
  assign T_4301 = T_4300 & T_1360_16;
  assign T_4304 = T_4271 & T_1365_17;
  assign T_4305 = T_4304 & T_1365_16;
  assign T_4308 = T_4275 & T_1370_17;
  assign T_4309 = T_4308 & T_1370_16;
  assign T_4312 = T_4279 & T_1375_17;
  assign T_4313 = T_4312 & T_1375_16;
  assign T_4315 = T_3830 & T_1360_18;
  assign T_4316 = T_4315 & T_1360_17;
  assign T_4317 = T_4316 & T_1360_16;
  assign T_4319 = T_3836 & T_1365_18;
  assign T_4320 = T_4319 & T_1365_17;
  assign T_4321 = T_4320 & T_1365_16;
  assign T_4323 = T_3840 & T_1370_18;
  assign T_4324 = T_4323 & T_1370_17;
  assign T_4325 = T_4324 & T_1370_16;
  assign T_4327 = T_3846 & T_1375_18;
  assign T_4328 = T_4327 & T_1375_17;
  assign T_4329 = T_4328 & T_1375_16;
  assign T_4331 = T_3730 & T_1360_21;
  assign T_4333 = T_3736 & T_1365_21;
  assign T_4335 = T_3740 & T_1370_21;
  assign T_4337 = T_3746 & T_1375_21;
  assign T_4339 = T_3730 & T_1360_20;
  assign T_4341 = T_3736 & T_1365_20;
  assign T_4343 = T_3740 & T_1370_20;
  assign T_4345 = T_3746 & T_1375_20;
  assign T_4347 = T_3890 & T_1360_24;
  assign T_4348 = T_4347 & T_1360_23;
  assign T_4350 = T_3896 & T_1365_24;
  assign T_4351 = T_4350 & T_1365_23;
  assign T_4353 = T_3900 & T_1370_24;
  assign T_4354 = T_4353 & T_1370_23;
  assign T_4356 = T_3906 & T_1375_24;
  assign T_4357 = T_4356 & T_1375_23;
  assign T_4360 = T_4347 & T_1360_22;
  assign T_4363 = T_4350 & T_1365_22;
  assign T_4366 = T_4353 & T_1370_22;
  assign T_4369 = T_4356 & T_1375_22;
  assign T_4371 = T_3890 & T_1360_23;
  assign T_4372 = T_4371 & T_1360_22;
  assign T_4374 = T_3896 & T_1365_23;
  assign T_4375 = T_4374 & T_1365_22;
  assign T_4377 = T_3900 & T_1370_23;
  assign T_4378 = T_4377 & T_1370_22;
  assign T_4380 = T_3906 & T_1375_23;
  assign T_4381 = T_4380 & T_1375_22;
  assign T_4422_0 = T_1225;
  assign T_4422_1 = T_1270;
  assign T_4422_2 = 1'h1;
  assign T_4422_3 = 1'h1;
  assign T_4422_4 = T_1342;
  assign T_4422_5 = T_1234;
  assign T_4422_6 = T_1279;
  assign T_4422_7 = 1'h1;
  assign T_4422_8 = 1'h1;
  assign T_4422_9 = 1'h1;
  assign T_4422_10 = T_1243;
  assign T_4422_11 = T_1324;
  assign T_4422_12 = 1'h1;
  assign T_4422_13 = 1'h1;
  assign T_4422_14 = 1'h1;
  assign T_4422_15 = 1'h1;
  assign T_4422_16 = T_1315;
  assign T_4422_17 = 1'h1;
  assign T_4422_18 = T_1306;
  assign T_4422_19 = T_1333;
  assign T_4422_20 = T_1252;
  assign T_4422_21 = T_1297;
  assign T_4422_22 = 1'h1;
  assign T_4422_23 = 1'h1;
  assign T_4422_24 = 1'h1;
  assign T_4422_25 = 1'h1;
  assign T_4422_26 = 1'h1;
  assign T_4422_27 = 1'h1;
  assign T_4422_28 = T_1288;
  assign T_4422_29 = T_1261;
  assign T_4422_30 = 1'h1;
  assign T_4422_31 = 1'h1;
  assign T_4493_0 = {{20'd0}, ctrl_sck_div};
  assign T_4493_1 = {{30'd0}, T_1952};
  assign T_4493_2 = 32'h0;
  assign T_4493_3 = 32'h0;
  assign T_4493_4 = {{31'd0}, ctrl_cs_id};
  assign T_4493_5 = {{31'd0}, ctrl_cs_dflt_0};
  assign T_4493_6 = {{30'd0}, ctrl_cs_mode};
  assign T_4493_7 = 32'h0;
  assign T_4493_8 = 32'h0;
  assign T_4493_9 = 32'h0;
  assign T_4493_10 = {{8'd0}, T_1752};
  assign T_4493_11 = {{8'd0}, T_2472};
  assign T_4493_12 = 32'h0;
  assign T_4493_13 = 32'h0;
  assign T_4493_14 = 32'h0;
  assign T_4493_15 = 32'h0;
  assign T_4493_16 = {{12'd0}, T_2392};
  assign T_4493_17 = 32'h0;
  assign T_4493_18 = T_2228;
  assign T_4493_19 = T_2592;
  assign T_4493_20 = {{28'd0}, ctrl_wm_tx};
  assign T_4493_21 = {{28'd0}, ctrl_wm_rx};
  assign T_4493_22 = 32'h0;
  assign T_4493_23 = 32'h0;
  assign T_4493_24 = 32'h0;
  assign T_4493_25 = 32'h0;
  assign T_4493_26 = 32'h0;
  assign T_4493_27 = 32'h0;
  assign T_4493_28 = {{30'd0}, T_2072};
  assign T_4493_29 = {{30'd0}, T_1872};
  assign T_4493_30 = 32'h0;
  assign T_4493_31 = 32'h0;
  assign GEN_4 = GEN_178;
  assign GEN_148 = 5'h1 == T_3414 ? T_4422_1 : T_4422_0;
  assign GEN_149 = 5'h2 == T_3414 ? T_4422_2 : GEN_148;
  assign GEN_150 = 5'h3 == T_3414 ? T_4422_3 : GEN_149;
  assign GEN_151 = 5'h4 == T_3414 ? T_4422_4 : GEN_150;
  assign GEN_152 = 5'h5 == T_3414 ? T_4422_5 : GEN_151;
  assign GEN_153 = 5'h6 == T_3414 ? T_4422_6 : GEN_152;
  assign GEN_154 = 5'h7 == T_3414 ? T_4422_7 : GEN_153;
  assign GEN_155 = 5'h8 == T_3414 ? T_4422_8 : GEN_154;
  assign GEN_156 = 5'h9 == T_3414 ? T_4422_9 : GEN_155;
  assign GEN_157 = 5'ha == T_3414 ? T_4422_10 : GEN_156;
  assign GEN_158 = 5'hb == T_3414 ? T_4422_11 : GEN_157;
  assign GEN_159 = 5'hc == T_3414 ? T_4422_12 : GEN_158;
  assign GEN_160 = 5'hd == T_3414 ? T_4422_13 : GEN_159;
  assign GEN_161 = 5'he == T_3414 ? T_4422_14 : GEN_160;
  assign GEN_162 = 5'hf == T_3414 ? T_4422_15 : GEN_161;
  assign GEN_163 = 5'h10 == T_3414 ? T_4422_16 : GEN_162;
  assign GEN_164 = 5'h11 == T_3414 ? T_4422_17 : GEN_163;
  assign GEN_165 = 5'h12 == T_3414 ? T_4422_18 : GEN_164;
  assign GEN_166 = 5'h13 == T_3414 ? T_4422_19 : GEN_165;
  assign GEN_167 = 5'h14 == T_3414 ? T_4422_20 : GEN_166;
  assign GEN_168 = 5'h15 == T_3414 ? T_4422_21 : GEN_167;
  assign GEN_169 = 5'h16 == T_3414 ? T_4422_22 : GEN_168;
  assign GEN_170 = 5'h17 == T_3414 ? T_4422_23 : GEN_169;
  assign GEN_171 = 5'h18 == T_3414 ? T_4422_24 : GEN_170;
  assign GEN_172 = 5'h19 == T_3414 ? T_4422_25 : GEN_171;
  assign GEN_173 = 5'h1a == T_3414 ? T_4422_26 : GEN_172;
  assign GEN_174 = 5'h1b == T_3414 ? T_4422_27 : GEN_173;
  assign GEN_175 = 5'h1c == T_3414 ? T_4422_28 : GEN_174;
  assign GEN_176 = 5'h1d == T_3414 ? T_4422_29 : GEN_175;
  assign GEN_177 = 5'h1e == T_3414 ? T_4422_30 : GEN_176;
  assign GEN_178 = 5'h1f == T_3414 ? T_4422_31 : GEN_177;
  assign GEN_5 = GEN_209;
  assign GEN_179 = 5'h1 == T_3414 ? T_4493_1 : T_4493_0;
  assign GEN_180 = 5'h2 == T_3414 ? T_4493_2 : GEN_179;
  assign GEN_181 = 5'h3 == T_3414 ? T_4493_3 : GEN_180;
  assign GEN_182 = 5'h4 == T_3414 ? T_4493_4 : GEN_181;
  assign GEN_183 = 5'h5 == T_3414 ? T_4493_5 : GEN_182;
  assign GEN_184 = 5'h6 == T_3414 ? T_4493_6 : GEN_183;
  assign GEN_185 = 5'h7 == T_3414 ? T_4493_7 : GEN_184;
  assign GEN_186 = 5'h8 == T_3414 ? T_4493_8 : GEN_185;
  assign GEN_187 = 5'h9 == T_3414 ? T_4493_9 : GEN_186;
  assign GEN_188 = 5'ha == T_3414 ? T_4493_10 : GEN_187;
  assign GEN_189 = 5'hb == T_3414 ? T_4493_11 : GEN_188;
  assign GEN_190 = 5'hc == T_3414 ? T_4493_12 : GEN_189;
  assign GEN_191 = 5'hd == T_3414 ? T_4493_13 : GEN_190;
  assign GEN_192 = 5'he == T_3414 ? T_4493_14 : GEN_191;
  assign GEN_193 = 5'hf == T_3414 ? T_4493_15 : GEN_192;
  assign GEN_194 = 5'h10 == T_3414 ? T_4493_16 : GEN_193;
  assign GEN_195 = 5'h11 == T_3414 ? T_4493_17 : GEN_194;
  assign GEN_196 = 5'h12 == T_3414 ? T_4493_18 : GEN_195;
  assign GEN_197 = 5'h13 == T_3414 ? T_4493_19 : GEN_196;
  assign GEN_198 = 5'h14 == T_3414 ? T_4493_20 : GEN_197;
  assign GEN_199 = 5'h15 == T_3414 ? T_4493_21 : GEN_198;
  assign GEN_200 = 5'h16 == T_3414 ? T_4493_22 : GEN_199;
  assign GEN_201 = 5'h17 == T_3414 ? T_4493_23 : GEN_200;
  assign GEN_202 = 5'h18 == T_3414 ? T_4493_24 : GEN_201;
  assign GEN_203 = 5'h19 == T_3414 ? T_4493_25 : GEN_202;
  assign GEN_204 = 5'h1a == T_3414 ? T_4493_26 : GEN_203;
  assign GEN_205 = 5'h1b == T_3414 ? T_4493_27 : GEN_204;
  assign GEN_206 = 5'h1c == T_3414 ? T_4493_28 : GEN_205;
  assign GEN_207 = 5'h1d == T_3414 ? T_4493_29 : GEN_206;
  assign GEN_208 = 5'h1e == T_3414 ? T_4493_30 : GEN_207;
  assign GEN_209 = 5'h1f == T_3414 ? T_4493_31 : GEN_208;
  assign T_4530 = GEN_4 ? GEN_5 : 32'h0;
  assign T_4531 = T_1102_bits_extra[9:8];
  assign T_4533 = T_1102_bits_extra[7:3];
  assign T_4534 = T_1102_bits_extra[2:0];
  assign T_4545_opcode = 3'h0;
  assign T_4545_param = 2'h0;
  assign T_4545_size = T_4534;
  assign T_4545_source = T_4533;
  assign T_4545_sink = 1'h0;
  assign T_4545_addr_lo = T_4531;
  assign T_4545_data = 32'h0;
  assign T_4545_error = 1'h0;

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_fmt_proto <= T_955_fmt_proto;
    end else begin
      if (T_2252) begin
        ctrl_fmt_proto <= T_1973;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_fmt_endian <= T_955_fmt_endian;
    end else begin
      if (T_2292) begin
        ctrl_fmt_endian <= T_2293;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_fmt_iodir <= T_955_fmt_iodir;
    end else begin
      if (T_2332) begin
        ctrl_fmt_iodir <= T_2333;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_fmt_len <= T_955_fmt_len;
    end else begin
      if (T_2372) begin
        ctrl_fmt_len <= T_2373;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_sck_div <= T_955_sck_div;
    end else begin
      if (T_1612) begin
        ctrl_sck_div <= T_1613;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_sck_pol <= T_955_sck_pol;
    end else begin
      if (T_1932) begin
        ctrl_sck_pol <= T_1853;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_sck_pha <= T_955_sck_pha;
    end else begin
      if (T_1892) begin
        ctrl_sck_pha <= T_1653;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_cs_id <= T_955_cs_id;
    end else begin
      if (T_2612) begin
        ctrl_cs_id <= T_1653;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_cs_dflt_0 <= T_955_cs_dflt_0;
    end else begin
      if (T_1652) begin
        ctrl_cs_dflt_0 <= T_1653;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_cs_mode <= T_955_cs_mode;
    end else begin
      if (T_1972) begin
        ctrl_cs_mode <= T_1973;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_dla_cssck <= T_955_dla_cssck;
    end else begin
      if (T_1692) begin
        ctrl_dla_cssck <= T_1693;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_dla_sckcs <= T_955_dla_sckcs;
    end else begin
      if (T_1732) begin
        ctrl_dla_sckcs <= T_1733;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_dla_intercs <= T_955_dla_intercs;
    end else begin
      if (T_2412) begin
        ctrl_dla_intercs <= T_1693;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_dla_interxfr <= T_955_dla_interxfr;
    end else begin
      if (T_2452) begin
        ctrl_dla_interxfr <= T_1733;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_wm_tx <= T_955_wm_tx;
    end else begin
      if (T_1772) begin
        ctrl_wm_tx <= T_1773;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_wm_rx <= T_955_wm_rx;
    end else begin
      if (T_2092) begin
        ctrl_wm_rx <= T_1773;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ie_txwm <= T_1021_txwm;
    end else begin
      if (T_2012) begin
        ie_txwm <= T_1653;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ie_rxwm <= T_1021_rxwm;
    end else begin
      if (T_2052) begin
        ie_rxwm <= T_1853;
      end
    end
endmodule
