 /*                                                                      
 Copyright 2017 Silicon Integrated Microelectronics, Inc.                
                                                                         
 Licensed under the Apache License, Version 2.0 (the "License");         
 you may not use this file except in compliance with the License.        
 You may obtain a copy of the License at                                 
                                                                         
     http://www.apache.org/licenses/LICENSE-2.0                          
                                                                         
  Unless required by applicable law or agreed to in writing, software    
 distributed under the License is distributed on an "AS IS" BASIS,       
 WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 See the License for the specific language governing permissions and     
 limitations under the License.                                          
 */                                                                      
                                                                         
                                                                         
                                                                         
module sirv_gpio(
  input   clock,
  input   reset,
  output  io_interrupts_0_0,
  output  io_interrupts_0_1,
  output  io_interrupts_0_2,
  output  io_interrupts_0_3,
  output  io_interrupts_0_4,
  output  io_interrupts_0_5,
  output  io_interrupts_0_6,
  output  io_interrupts_0_7,
  output  io_interrupts_0_8,
  output  io_interrupts_0_9,
  output  io_interrupts_0_10,
  output  io_interrupts_0_11,
  output  io_interrupts_0_12,
  output  io_interrupts_0_13,
  output  io_interrupts_0_14,
  output  io_interrupts_0_15,
  output  io_interrupts_0_16,
  output  io_interrupts_0_17,
  output  io_interrupts_0_18,
  output  io_interrupts_0_19,
  output  io_interrupts_0_20,
  output  io_interrupts_0_21,
  output  io_interrupts_0_22,
  output  io_interrupts_0_23,
  output  io_interrupts_0_24,
  output  io_interrupts_0_25,
  output  io_interrupts_0_26,
  output  io_interrupts_0_27,
  output  io_interrupts_0_28,
  output  io_interrupts_0_29,
  output  io_interrupts_0_30,
  output  io_interrupts_0_31,
  output  io_in_0_a_ready,
  input   io_in_0_a_valid,
  input  [2:0] io_in_0_a_bits_opcode,
  input  [2:0] io_in_0_a_bits_param,
  input  [2:0] io_in_0_a_bits_size,
  input  [4:0] io_in_0_a_bits_source,
  input  [28:0] io_in_0_a_bits_address,
  input  [3:0] io_in_0_a_bits_mask,
  input  [31:0] io_in_0_a_bits_data,
  input   io_in_0_b_ready,
  output  io_in_0_b_valid,
  output [2:0] io_in_0_b_bits_opcode,
  output [1:0] io_in_0_b_bits_param,
  output [2:0] io_in_0_b_bits_size,
  output [4:0] io_in_0_b_bits_source,
  output [28:0] io_in_0_b_bits_address,
  output [3:0] io_in_0_b_bits_mask,
  output [31:0] io_in_0_b_bits_data,
  output  io_in_0_c_ready,
  input   io_in_0_c_valid,
  input  [2:0] io_in_0_c_bits_opcode,
  input  [2:0] io_in_0_c_bits_param,
  input  [2:0] io_in_0_c_bits_size,
  input  [4:0] io_in_0_c_bits_source,
  input  [28:0] io_in_0_c_bits_address,
  input  [31:0] io_in_0_c_bits_data,
  input   io_in_0_c_bits_error,
  input   io_in_0_d_ready,
  output  io_in_0_d_valid,
  output [2:0] io_in_0_d_bits_opcode,
  output [1:0] io_in_0_d_bits_param,
  output [2:0] io_in_0_d_bits_size,
  output [4:0] io_in_0_d_bits_source,
  output  io_in_0_d_bits_sink,
  output [1:0] io_in_0_d_bits_addr_lo,
  output [31:0] io_in_0_d_bits_data,
  output  io_in_0_d_bits_error,
  output  io_in_0_e_ready,
  input   io_in_0_e_valid,
  input   io_in_0_e_bits_sink,
  input   io_port_pins_0_i_ival,
  output  io_port_pins_0_o_oval,
  output  io_port_pins_0_o_oe,
  output  io_port_pins_0_o_ie,
  output  io_port_pins_0_o_pue,
  output  io_port_pins_0_o_ds,
  input   io_port_pins_1_i_ival,
  output  io_port_pins_1_o_oval,
  output  io_port_pins_1_o_oe,
  output  io_port_pins_1_o_ie,
  output  io_port_pins_1_o_pue,
  output  io_port_pins_1_o_ds,
  input   io_port_pins_2_i_ival,
  output  io_port_pins_2_o_oval,
  output  io_port_pins_2_o_oe,
  output  io_port_pins_2_o_ie,
  output  io_port_pins_2_o_pue,
  output  io_port_pins_2_o_ds,
  input   io_port_pins_3_i_ival,
  output  io_port_pins_3_o_oval,
  output  io_port_pins_3_o_oe,
  output  io_port_pins_3_o_ie,
  output  io_port_pins_3_o_pue,
  output  io_port_pins_3_o_ds,
  input   io_port_pins_4_i_ival,
  output  io_port_pins_4_o_oval,
  output  io_port_pins_4_o_oe,
  output  io_port_pins_4_o_ie,
  output  io_port_pins_4_o_pue,
  output  io_port_pins_4_o_ds,
  input   io_port_pins_5_i_ival,
  output  io_port_pins_5_o_oval,
  output  io_port_pins_5_o_oe,
  output  io_port_pins_5_o_ie,
  output  io_port_pins_5_o_pue,
  output  io_port_pins_5_o_ds,
  input   io_port_pins_6_i_ival,
  output  io_port_pins_6_o_oval,
  output  io_port_pins_6_o_oe,
  output  io_port_pins_6_o_ie,
  output  io_port_pins_6_o_pue,
  output  io_port_pins_6_o_ds,
  input   io_port_pins_7_i_ival,
  output  io_port_pins_7_o_oval,
  output  io_port_pins_7_o_oe,
  output  io_port_pins_7_o_ie,
  output  io_port_pins_7_o_pue,
  output  io_port_pins_7_o_ds,
  input   io_port_pins_8_i_ival,
  output  io_port_pins_8_o_oval,
  output  io_port_pins_8_o_oe,
  output  io_port_pins_8_o_ie,
  output  io_port_pins_8_o_pue,
  output  io_port_pins_8_o_ds,
  input   io_port_pins_9_i_ival,
  output  io_port_pins_9_o_oval,
  output  io_port_pins_9_o_oe,
  output  io_port_pins_9_o_ie,
  output  io_port_pins_9_o_pue,
  output  io_port_pins_9_o_ds,
  input   io_port_pins_10_i_ival,
  output  io_port_pins_10_o_oval,
  output  io_port_pins_10_o_oe,
  output  io_port_pins_10_o_ie,
  output  io_port_pins_10_o_pue,
  output  io_port_pins_10_o_ds,
  input   io_port_pins_11_i_ival,
  output  io_port_pins_11_o_oval,
  output  io_port_pins_11_o_oe,
  output  io_port_pins_11_o_ie,
  output  io_port_pins_11_o_pue,
  output  io_port_pins_11_o_ds,
  input   io_port_pins_12_i_ival,
  output  io_port_pins_12_o_oval,
  output  io_port_pins_12_o_oe,
  output  io_port_pins_12_o_ie,
  output  io_port_pins_12_o_pue,
  output  io_port_pins_12_o_ds,
  input   io_port_pins_13_i_ival,
  output  io_port_pins_13_o_oval,
  output  io_port_pins_13_o_oe,
  output  io_port_pins_13_o_ie,
  output  io_port_pins_13_o_pue,
  output  io_port_pins_13_o_ds,
  input   io_port_pins_14_i_ival,
  output  io_port_pins_14_o_oval,
  output  io_port_pins_14_o_oe,
  output  io_port_pins_14_o_ie,
  output  io_port_pins_14_o_pue,
  output  io_port_pins_14_o_ds,
  input   io_port_pins_15_i_ival,
  output  io_port_pins_15_o_oval,
  output  io_port_pins_15_o_oe,
  output  io_port_pins_15_o_ie,
  output  io_port_pins_15_o_pue,
  output  io_port_pins_15_o_ds,
  input   io_port_pins_16_i_ival,
  output  io_port_pins_16_o_oval,
  output  io_port_pins_16_o_oe,
  output  io_port_pins_16_o_ie,
  output  io_port_pins_16_o_pue,
  output  io_port_pins_16_o_ds,
  input   io_port_pins_17_i_ival,
  output  io_port_pins_17_o_oval,
  output  io_port_pins_17_o_oe,
  output  io_port_pins_17_o_ie,
  output  io_port_pins_17_o_pue,
  output  io_port_pins_17_o_ds,
  input   io_port_pins_18_i_ival,
  output  io_port_pins_18_o_oval,
  output  io_port_pins_18_o_oe,
  output  io_port_pins_18_o_ie,
  output  io_port_pins_18_o_pue,
  output  io_port_pins_18_o_ds,
  input   io_port_pins_19_i_ival,
  output  io_port_pins_19_o_oval,
  output  io_port_pins_19_o_oe,
  output  io_port_pins_19_o_ie,
  output  io_port_pins_19_o_pue,
  output  io_port_pins_19_o_ds,
  input   io_port_pins_20_i_ival,
  output  io_port_pins_20_o_oval,
  output  io_port_pins_20_o_oe,
  output  io_port_pins_20_o_ie,
  output  io_port_pins_20_o_pue,
  output  io_port_pins_20_o_ds,
  input   io_port_pins_21_i_ival,
  output  io_port_pins_21_o_oval,
  output  io_port_pins_21_o_oe,
  output  io_port_pins_21_o_ie,
  output  io_port_pins_21_o_pue,
  output  io_port_pins_21_o_ds,
  input   io_port_pins_22_i_ival,
  output  io_port_pins_22_o_oval,
  output  io_port_pins_22_o_oe,
  output  io_port_pins_22_o_ie,
  output  io_port_pins_22_o_pue,
  output  io_port_pins_22_o_ds,
  input   io_port_pins_23_i_ival,
  output  io_port_pins_23_o_oval,
  output  io_port_pins_23_o_oe,
  output  io_port_pins_23_o_ie,
  output  io_port_pins_23_o_pue,
  output  io_port_pins_23_o_ds,
  input   io_port_pins_24_i_ival,
  output  io_port_pins_24_o_oval,
  output  io_port_pins_24_o_oe,
  output  io_port_pins_24_o_ie,
  output  io_port_pins_24_o_pue,
  output  io_port_pins_24_o_ds,
  input   io_port_pins_25_i_ival,
  output  io_port_pins_25_o_oval,
  output  io_port_pins_25_o_oe,
  output  io_port_pins_25_o_ie,
  output  io_port_pins_25_o_pue,
  output  io_port_pins_25_o_ds,
  input   io_port_pins_26_i_ival,
  output  io_port_pins_26_o_oval,
  output  io_port_pins_26_o_oe,
  output  io_port_pins_26_o_ie,
  output  io_port_pins_26_o_pue,
  output  io_port_pins_26_o_ds,
  input   io_port_pins_27_i_ival,
  output  io_port_pins_27_o_oval,
  output  io_port_pins_27_o_oe,
  output  io_port_pins_27_o_ie,
  output  io_port_pins_27_o_pue,
  output  io_port_pins_27_o_ds,
  input   io_port_pins_28_i_ival,
  output  io_port_pins_28_o_oval,
  output  io_port_pins_28_o_oe,
  output  io_port_pins_28_o_ie,
  output  io_port_pins_28_o_pue,
  output  io_port_pins_28_o_ds,
  input   io_port_pins_29_i_ival,
  output  io_port_pins_29_o_oval,
  output  io_port_pins_29_o_oe,
  output  io_port_pins_29_o_ie,
  output  io_port_pins_29_o_pue,
  output  io_port_pins_29_o_ds,
  input   io_port_pins_30_i_ival,
  output  io_port_pins_30_o_oval,
  output  io_port_pins_30_o_oe,
  output  io_port_pins_30_o_ie,
  output  io_port_pins_30_o_pue,
  output  io_port_pins_30_o_ds,
  input   io_port_pins_31_i_ival,
  output  io_port_pins_31_o_oval,
  output  io_port_pins_31_o_oe,
  output  io_port_pins_31_o_ie,
  output  io_port_pins_31_o_pue,
  output  io_port_pins_31_o_ds,
  output  io_port_iof_0_0_i_ival,
  input   io_port_iof_0_0_o_oval,
  input   io_port_iof_0_0_o_oe,
  input   io_port_iof_0_0_o_ie,
  input   io_port_iof_0_0_o_valid,
  output  io_port_iof_0_1_i_ival,
  input   io_port_iof_0_1_o_oval,
  input   io_port_iof_0_1_o_oe,
  input   io_port_iof_0_1_o_ie,
  input   io_port_iof_0_1_o_valid,
  output  io_port_iof_0_2_i_ival,
  input   io_port_iof_0_2_o_oval,
  input   io_port_iof_0_2_o_oe,
  input   io_port_iof_0_2_o_ie,
  input   io_port_iof_0_2_o_valid,
  output  io_port_iof_0_3_i_ival,
  input   io_port_iof_0_3_o_oval,
  input   io_port_iof_0_3_o_oe,
  input   io_port_iof_0_3_o_ie,
  input   io_port_iof_0_3_o_valid,
  output  io_port_iof_0_4_i_ival,
  input   io_port_iof_0_4_o_oval,
  input   io_port_iof_0_4_o_oe,
  input   io_port_iof_0_4_o_ie,
  input   io_port_iof_0_4_o_valid,
  output  io_port_iof_0_5_i_ival,
  input   io_port_iof_0_5_o_oval,
  input   io_port_iof_0_5_o_oe,
  input   io_port_iof_0_5_o_ie,
  input   io_port_iof_0_5_o_valid,
  output  io_port_iof_0_6_i_ival,
  input   io_port_iof_0_6_o_oval,
  input   io_port_iof_0_6_o_oe,
  input   io_port_iof_0_6_o_ie,
  input   io_port_iof_0_6_o_valid,
  output  io_port_iof_0_7_i_ival,
  input   io_port_iof_0_7_o_oval,
  input   io_port_iof_0_7_o_oe,
  input   io_port_iof_0_7_o_ie,
  input   io_port_iof_0_7_o_valid,
  output  io_port_iof_0_8_i_ival,
  input   io_port_iof_0_8_o_oval,
  input   io_port_iof_0_8_o_oe,
  input   io_port_iof_0_8_o_ie,
  input   io_port_iof_0_8_o_valid,
  output  io_port_iof_0_9_i_ival,
  input   io_port_iof_0_9_o_oval,
  input   io_port_iof_0_9_o_oe,
  input   io_port_iof_0_9_o_ie,
  input   io_port_iof_0_9_o_valid,
  output  io_port_iof_0_10_i_ival,
  input   io_port_iof_0_10_o_oval,
  input   io_port_iof_0_10_o_oe,
  input   io_port_iof_0_10_o_ie,
  input   io_port_iof_0_10_o_valid,
  output  io_port_iof_0_11_i_ival,
  input   io_port_iof_0_11_o_oval,
  input   io_port_iof_0_11_o_oe,
  input   io_port_iof_0_11_o_ie,
  input   io_port_iof_0_11_o_valid,
  output  io_port_iof_0_12_i_ival,
  input   io_port_iof_0_12_o_oval,
  input   io_port_iof_0_12_o_oe,
  input   io_port_iof_0_12_o_ie,
  input   io_port_iof_0_12_o_valid,
  output  io_port_iof_0_13_i_ival,
  input   io_port_iof_0_13_o_oval,
  input   io_port_iof_0_13_o_oe,
  input   io_port_iof_0_13_o_ie,
  input   io_port_iof_0_13_o_valid,
  output  io_port_iof_0_14_i_ival,
  input   io_port_iof_0_14_o_oval,
  input   io_port_iof_0_14_o_oe,
  input   io_port_iof_0_14_o_ie,
  input   io_port_iof_0_14_o_valid,
  output  io_port_iof_0_15_i_ival,
  input   io_port_iof_0_15_o_oval,
  input   io_port_iof_0_15_o_oe,
  input   io_port_iof_0_15_o_ie,
  input   io_port_iof_0_15_o_valid,
  output  io_port_iof_0_16_i_ival,
  input   io_port_iof_0_16_o_oval,
  input   io_port_iof_0_16_o_oe,
  input   io_port_iof_0_16_o_ie,
  input   io_port_iof_0_16_o_valid,
  output  io_port_iof_0_17_i_ival,
  input   io_port_iof_0_17_o_oval,
  input   io_port_iof_0_17_o_oe,
  input   io_port_iof_0_17_o_ie,
  input   io_port_iof_0_17_o_valid,
  output  io_port_iof_0_18_i_ival,
  input   io_port_iof_0_18_o_oval,
  input   io_port_iof_0_18_o_oe,
  input   io_port_iof_0_18_o_ie,
  input   io_port_iof_0_18_o_valid,
  output  io_port_iof_0_19_i_ival,
  input   io_port_iof_0_19_o_oval,
  input   io_port_iof_0_19_o_oe,
  input   io_port_iof_0_19_o_ie,
  input   io_port_iof_0_19_o_valid,
  output  io_port_iof_0_20_i_ival,
  input   io_port_iof_0_20_o_oval,
  input   io_port_iof_0_20_o_oe,
  input   io_port_iof_0_20_o_ie,
  input   io_port_iof_0_20_o_valid,
  output  io_port_iof_0_21_i_ival,
  input   io_port_iof_0_21_o_oval,
  input   io_port_iof_0_21_o_oe,
  input   io_port_iof_0_21_o_ie,
  input   io_port_iof_0_21_o_valid,
  output  io_port_iof_0_22_i_ival,
  input   io_port_iof_0_22_o_oval,
  input   io_port_iof_0_22_o_oe,
  input   io_port_iof_0_22_o_ie,
  input   io_port_iof_0_22_o_valid,
  output  io_port_iof_0_23_i_ival,
  input   io_port_iof_0_23_o_oval,
  input   io_port_iof_0_23_o_oe,
  input   io_port_iof_0_23_o_ie,
  input   io_port_iof_0_23_o_valid,
  output  io_port_iof_0_24_i_ival,
  input   io_port_iof_0_24_o_oval,
  input   io_port_iof_0_24_o_oe,
  input   io_port_iof_0_24_o_ie,
  input   io_port_iof_0_24_o_valid,
  output  io_port_iof_0_25_i_ival,
  input   io_port_iof_0_25_o_oval,
  input   io_port_iof_0_25_o_oe,
  input   io_port_iof_0_25_o_ie,
  input   io_port_iof_0_25_o_valid,
  output  io_port_iof_0_26_i_ival,
  input   io_port_iof_0_26_o_oval,
  input   io_port_iof_0_26_o_oe,
  input   io_port_iof_0_26_o_ie,
  input   io_port_iof_0_26_o_valid,
  output  io_port_iof_0_27_i_ival,
  input   io_port_iof_0_27_o_oval,
  input   io_port_iof_0_27_o_oe,
  input   io_port_iof_0_27_o_ie,
  input   io_port_iof_0_27_o_valid,
  output  io_port_iof_0_28_i_ival,
  input   io_port_iof_0_28_o_oval,
  input   io_port_iof_0_28_o_oe,
  input   io_port_iof_0_28_o_ie,
  input   io_port_iof_0_28_o_valid,
  output  io_port_iof_0_29_i_ival,
  input   io_port_iof_0_29_o_oval,
  input   io_port_iof_0_29_o_oe,
  input   io_port_iof_0_29_o_ie,
  input   io_port_iof_0_29_o_valid,
  output  io_port_iof_0_30_i_ival,
  input   io_port_iof_0_30_o_oval,
  input   io_port_iof_0_30_o_oe,
  input   io_port_iof_0_30_o_ie,
  input   io_port_iof_0_30_o_valid,
  output  io_port_iof_0_31_i_ival,
  input   io_port_iof_0_31_o_oval,
  input   io_port_iof_0_31_o_oe,
  input   io_port_iof_0_31_o_ie,
  input   io_port_iof_0_31_o_valid,
  output  io_port_iof_1_0_i_ival,
  input   io_port_iof_1_0_o_oval,
  input   io_port_iof_1_0_o_oe,
  input   io_port_iof_1_0_o_ie,
  input   io_port_iof_1_0_o_valid,
  output  io_port_iof_1_1_i_ival,
  input   io_port_iof_1_1_o_oval,
  input   io_port_iof_1_1_o_oe,
  input   io_port_iof_1_1_o_ie,
  input   io_port_iof_1_1_o_valid,
  output  io_port_iof_1_2_i_ival,
  input   io_port_iof_1_2_o_oval,
  input   io_port_iof_1_2_o_oe,
  input   io_port_iof_1_2_o_ie,
  input   io_port_iof_1_2_o_valid,
  output  io_port_iof_1_3_i_ival,
  input   io_port_iof_1_3_o_oval,
  input   io_port_iof_1_3_o_oe,
  input   io_port_iof_1_3_o_ie,
  input   io_port_iof_1_3_o_valid,
  output  io_port_iof_1_4_i_ival,
  input   io_port_iof_1_4_o_oval,
  input   io_port_iof_1_4_o_oe,
  input   io_port_iof_1_4_o_ie,
  input   io_port_iof_1_4_o_valid,
  output  io_port_iof_1_5_i_ival,
  input   io_port_iof_1_5_o_oval,
  input   io_port_iof_1_5_o_oe,
  input   io_port_iof_1_5_o_ie,
  input   io_port_iof_1_5_o_valid,
  output  io_port_iof_1_6_i_ival,
  input   io_port_iof_1_6_o_oval,
  input   io_port_iof_1_6_o_oe,
  input   io_port_iof_1_6_o_ie,
  input   io_port_iof_1_6_o_valid,
  output  io_port_iof_1_7_i_ival,
  input   io_port_iof_1_7_o_oval,
  input   io_port_iof_1_7_o_oe,
  input   io_port_iof_1_7_o_ie,
  input   io_port_iof_1_7_o_valid,
  output  io_port_iof_1_8_i_ival,
  input   io_port_iof_1_8_o_oval,
  input   io_port_iof_1_8_o_oe,
  input   io_port_iof_1_8_o_ie,
  input   io_port_iof_1_8_o_valid,
  output  io_port_iof_1_9_i_ival,
  input   io_port_iof_1_9_o_oval,
  input   io_port_iof_1_9_o_oe,
  input   io_port_iof_1_9_o_ie,
  input   io_port_iof_1_9_o_valid,
  output  io_port_iof_1_10_i_ival,
  input   io_port_iof_1_10_o_oval,
  input   io_port_iof_1_10_o_oe,
  input   io_port_iof_1_10_o_ie,
  input   io_port_iof_1_10_o_valid,
  output  io_port_iof_1_11_i_ival,
  input   io_port_iof_1_11_o_oval,
  input   io_port_iof_1_11_o_oe,
  input   io_port_iof_1_11_o_ie,
  input   io_port_iof_1_11_o_valid,
  output  io_port_iof_1_12_i_ival,
  input   io_port_iof_1_12_o_oval,
  input   io_port_iof_1_12_o_oe,
  input   io_port_iof_1_12_o_ie,
  input   io_port_iof_1_12_o_valid,
  output  io_port_iof_1_13_i_ival,
  input   io_port_iof_1_13_o_oval,
  input   io_port_iof_1_13_o_oe,
  input   io_port_iof_1_13_o_ie,
  input   io_port_iof_1_13_o_valid,
  output  io_port_iof_1_14_i_ival,
  input   io_port_iof_1_14_o_oval,
  input   io_port_iof_1_14_o_oe,
  input   io_port_iof_1_14_o_ie,
  input   io_port_iof_1_14_o_valid,
  output  io_port_iof_1_15_i_ival,
  input   io_port_iof_1_15_o_oval,
  input   io_port_iof_1_15_o_oe,
  input   io_port_iof_1_15_o_ie,
  input   io_port_iof_1_15_o_valid,
  output  io_port_iof_1_16_i_ival,
  input   io_port_iof_1_16_o_oval,
  input   io_port_iof_1_16_o_oe,
  input   io_port_iof_1_16_o_ie,
  input   io_port_iof_1_16_o_valid,
  output  io_port_iof_1_17_i_ival,
  input   io_port_iof_1_17_o_oval,
  input   io_port_iof_1_17_o_oe,
  input   io_port_iof_1_17_o_ie,
  input   io_port_iof_1_17_o_valid,
  output  io_port_iof_1_18_i_ival,
  input   io_port_iof_1_18_o_oval,
  input   io_port_iof_1_18_o_oe,
  input   io_port_iof_1_18_o_ie,
  input   io_port_iof_1_18_o_valid,
  output  io_port_iof_1_19_i_ival,
  input   io_port_iof_1_19_o_oval,
  input   io_port_iof_1_19_o_oe,
  input   io_port_iof_1_19_o_ie,
  input   io_port_iof_1_19_o_valid,
  output  io_port_iof_1_20_i_ival,
  input   io_port_iof_1_20_o_oval,
  input   io_port_iof_1_20_o_oe,
  input   io_port_iof_1_20_o_ie,
  input   io_port_iof_1_20_o_valid,
  output  io_port_iof_1_21_i_ival,
  input   io_port_iof_1_21_o_oval,
  input   io_port_iof_1_21_o_oe,
  input   io_port_iof_1_21_o_ie,
  input   io_port_iof_1_21_o_valid,
  output  io_port_iof_1_22_i_ival,
  input   io_port_iof_1_22_o_oval,
  input   io_port_iof_1_22_o_oe,
  input   io_port_iof_1_22_o_ie,
  input   io_port_iof_1_22_o_valid,
  output  io_port_iof_1_23_i_ival,
  input   io_port_iof_1_23_o_oval,
  input   io_port_iof_1_23_o_oe,
  input   io_port_iof_1_23_o_ie,
  input   io_port_iof_1_23_o_valid,
  output  io_port_iof_1_24_i_ival,
  input   io_port_iof_1_24_o_oval,
  input   io_port_iof_1_24_o_oe,
  input   io_port_iof_1_24_o_ie,
  input   io_port_iof_1_24_o_valid,
  output  io_port_iof_1_25_i_ival,
  input   io_port_iof_1_25_o_oval,
  input   io_port_iof_1_25_o_oe,
  input   io_port_iof_1_25_o_ie,
  input   io_port_iof_1_25_o_valid,
  output  io_port_iof_1_26_i_ival,
  input   io_port_iof_1_26_o_oval,
  input   io_port_iof_1_26_o_oe,
  input   io_port_iof_1_26_o_ie,
  input   io_port_iof_1_26_o_valid,
  output  io_port_iof_1_27_i_ival,
  input   io_port_iof_1_27_o_oval,
  input   io_port_iof_1_27_o_oe,
  input   io_port_iof_1_27_o_ie,
  input   io_port_iof_1_27_o_valid,
  output  io_port_iof_1_28_i_ival,
  input   io_port_iof_1_28_o_oval,
  input   io_port_iof_1_28_o_oe,
  input   io_port_iof_1_28_o_ie,
  input   io_port_iof_1_28_o_valid,
  output  io_port_iof_1_29_i_ival,
  input   io_port_iof_1_29_o_oval,
  input   io_port_iof_1_29_o_oe,
  input   io_port_iof_1_29_o_ie,
  input   io_port_iof_1_29_o_valid,
  output  io_port_iof_1_30_i_ival,
  input   io_port_iof_1_30_o_oval,
  input   io_port_iof_1_30_o_oe,
  input   io_port_iof_1_30_o_ie,
  input   io_port_iof_1_30_o_valid,
  output  io_port_iof_1_31_i_ival,
  input   io_port_iof_1_31_o_oval,
  input   io_port_iof_1_31_o_oe,
  input   io_port_iof_1_31_o_ie,
  input   io_port_iof_1_31_o_valid
);
  reg [31:0] portReg;
  reg [31:0] GEN_399;
  wire  oeReg_clock;
  wire  oeReg_reset;
  wire [31:0] oeReg_io_d;
  wire [31:0] oeReg_io_q;
  wire  oeReg_io_en;
  wire  pueReg_clock;
  wire  pueReg_reset;
  wire [31:0] pueReg_io_d;
  wire [31:0] pueReg_io_q;
  wire  pueReg_io_en;
  reg [31:0] dsReg;
  reg [31:0] GEN_400;
  wire  ieReg_clock;
  wire  ieReg_reset;
  wire [31:0] ieReg_io_d;
  wire [31:0] ieReg_io_q;
  wire  ieReg_io_en;
  wire [31:0] inVal;
  wire  T_3188_0;
  wire  T_3188_1;
  wire  T_3188_2;
  wire  T_3188_3;
  wire  T_3188_4;
  wire  T_3188_5;
  wire  T_3188_6;
  wire  T_3188_7;
  wire  T_3188_8;
  wire  T_3188_9;
  wire  T_3188_10;
  wire  T_3188_11;
  wire  T_3188_12;
  wire  T_3188_13;
  wire  T_3188_14;
  wire  T_3188_15;
  wire  T_3188_16;
  wire  T_3188_17;
  wire  T_3188_18;
  wire  T_3188_19;
  wire  T_3188_20;
  wire  T_3188_21;
  wire  T_3188_22;
  wire  T_3188_23;
  wire  T_3188_24;
  wire  T_3188_25;
  wire  T_3188_26;
  wire  T_3188_27;
  wire  T_3188_28;
  wire  T_3188_29;
  wire  T_3188_30;
  wire  T_3188_31;
  wire [1:0] T_3223;
  wire [1:0] T_3224;
  wire [3:0] T_3225;
  wire [1:0] T_3226;
  wire [1:0] T_3227;
  wire [3:0] T_3228;
  wire [7:0] T_3229;
  wire [1:0] T_3230;
  wire [1:0] T_3231;
  wire [3:0] T_3232;
  wire [1:0] T_3233;
  wire [1:0] T_3234;
  wire [3:0] T_3235;
  wire [7:0] T_3236;
  wire [15:0] T_3237;
  wire [1:0] T_3238;
  wire [1:0] T_3239;
  wire [3:0] T_3240;
  wire [1:0] T_3241;
  wire [1:0] T_3242;
  wire [3:0] T_3243;
  wire [7:0] T_3244;
  wire [1:0] T_3245;
  wire [1:0] T_3246;
  wire [3:0] T_3247;
  wire [1:0] T_3248;
  wire [1:0] T_3249;
  wire [3:0] T_3250;
  wire [7:0] T_3251;
  wire [15:0] T_3252;
  wire [31:0] T_3253;
  reg [31:0] T_3256;
  reg [31:0] GEN_401;
  reg [31:0] T_3257;
  reg [31:0] GEN_402;
  reg [31:0] inSyncReg;
  reg [31:0] GEN_403;
  reg [31:0] valueReg;
  reg [31:0] GEN_404;
  reg [31:0] highIeReg;
  reg [31:0] GEN_405;
  reg [31:0] lowIeReg;
  reg [31:0] GEN_406;
  reg [31:0] riseIeReg;
  reg [31:0] GEN_407;
  reg [31:0] fallIeReg;
  reg [31:0] GEN_408;
  reg [31:0] highIpReg;
  reg [31:0] GEN_409;
  reg [31:0] lowIpReg;
  reg [31:0] GEN_410;
  reg [31:0] riseIpReg;
  reg [31:0] GEN_411;
  reg [31:0] fallIpReg;
  reg [31:0] GEN_412;
  wire  iofEnReg_clock;
  wire  iofEnReg_reset;
  wire [31:0] iofEnReg_io_d;
  wire [31:0] iofEnReg_io_q;
  wire  iofEnReg_io_en;
  reg [31:0] iofSelReg;
  reg [31:0] GEN_413;
  reg [31:0] xorReg;
  reg [31:0] GEN_414;
  wire [31:0] T_3269;
  wire [31:0] rise;
  wire [31:0] T_3270;
  wire [31:0] fall;
  wire  T_3295_ready;
  wire  T_3295_valid;
  wire  T_3295_bits_read;
  wire [9:0] T_3295_bits_index;
  wire [31:0] T_3295_bits_data;
  wire [3:0] T_3295_bits_mask;
  wire [9:0] T_3295_bits_extra;
  wire  T_3312;
  wire [26:0] T_3313;
  wire [1:0] T_3314;
  wire [6:0] T_3315;
  wire [9:0] T_3316;
  wire  T_3334_ready;
  wire  T_3334_valid;
  wire  T_3334_bits_read;
  wire [31:0] T_3334_bits_data;
  wire [9:0] T_3334_bits_extra;
  wire  T_3370_ready;
  wire  T_3370_valid;
  wire  T_3370_bits_read;
  wire [9:0] T_3370_bits_index;
  wire [31:0] T_3370_bits_data;
  wire [3:0] T_3370_bits_mask;
  wire [9:0] T_3370_bits_extra;
  wire [9:0] T_3455;
  wire  T_3457;
  wire [9:0] T_3463;
  wire [9:0] T_3464;
  wire  T_3466;
  wire [9:0] T_3472;
  wire [9:0] T_3473;
  wire  T_3475;
  wire [9:0] T_3481;
  wire [9:0] T_3482;
  wire  T_3484;
  wire [9:0] T_3490;
  wire [9:0] T_3491;
  wire  T_3493;
  wire [9:0] T_3499;
  wire [9:0] T_3500;
  wire  T_3502;
  wire [9:0] T_3508;
  wire [9:0] T_3509;
  wire  T_3511;
  wire [9:0] T_3517;
  wire [9:0] T_3518;
  wire  T_3520;
  wire [9:0] T_3526;
  wire [9:0] T_3527;
  wire  T_3529;
  wire [9:0] T_3535;
  wire [9:0] T_3536;
  wire  T_3538;
  wire [9:0] T_3544;
  wire [9:0] T_3545;
  wire  T_3547;
  wire [9:0] T_3553;
  wire [9:0] T_3554;
  wire  T_3556;
  wire [9:0] T_3562;
  wire [9:0] T_3563;
  wire  T_3565;
  wire [9:0] T_3571;
  wire [9:0] T_3572;
  wire  T_3574;
  wire [9:0] T_3580;
  wire [9:0] T_3581;
  wire  T_3583;
  wire [9:0] T_3589;
  wire [9:0] T_3590;
  wire  T_3592;
  wire [9:0] T_3598;
  wire [9:0] T_3599;
  wire  T_3601;
  wire  T_3609_0;
  wire  T_3609_1;
  wire  T_3609_2;
  wire  T_3609_3;
  wire  T_3609_4;
  wire  T_3609_5;
  wire  T_3609_6;
  wire  T_3609_7;
  wire  T_3609_8;
  wire  T_3609_9;
  wire  T_3609_10;
  wire  T_3609_11;
  wire  T_3609_12;
  wire  T_3609_13;
  wire  T_3609_14;
  wire  T_3609_15;
  wire  T_3609_16;
  wire  T_3614_0;
  wire  T_3614_1;
  wire  T_3614_2;
  wire  T_3614_3;
  wire  T_3614_4;
  wire  T_3614_5;
  wire  T_3614_6;
  wire  T_3614_7;
  wire  T_3614_8;
  wire  T_3614_9;
  wire  T_3614_10;
  wire  T_3614_11;
  wire  T_3614_12;
  wire  T_3614_13;
  wire  T_3614_14;
  wire  T_3614_15;
  wire  T_3614_16;
  wire  T_3619_0;
  wire  T_3619_1;
  wire  T_3619_2;
  wire  T_3619_3;
  wire  T_3619_4;
  wire  T_3619_5;
  wire  T_3619_6;
  wire  T_3619_7;
  wire  T_3619_8;
  wire  T_3619_9;
  wire  T_3619_10;
  wire  T_3619_11;
  wire  T_3619_12;
  wire  T_3619_13;
  wire  T_3619_14;
  wire  T_3619_15;
  wire  T_3619_16;
  wire  T_3624_0;
  wire  T_3624_1;
  wire  T_3624_2;
  wire  T_3624_3;
  wire  T_3624_4;
  wire  T_3624_5;
  wire  T_3624_6;
  wire  T_3624_7;
  wire  T_3624_8;
  wire  T_3624_9;
  wire  T_3624_10;
  wire  T_3624_11;
  wire  T_3624_12;
  wire  T_3624_13;
  wire  T_3624_14;
  wire  T_3624_15;
  wire  T_3624_16;
  wire  T_3629_0;
  wire  T_3629_1;
  wire  T_3629_2;
  wire  T_3629_3;
  wire  T_3629_4;
  wire  T_3629_5;
  wire  T_3629_6;
  wire  T_3629_7;
  wire  T_3629_8;
  wire  T_3629_9;
  wire  T_3629_10;
  wire  T_3629_11;
  wire  T_3629_12;
  wire  T_3629_13;
  wire  T_3629_14;
  wire  T_3629_15;
  wire  T_3629_16;
  wire  T_3634_0;
  wire  T_3634_1;
  wire  T_3634_2;
  wire  T_3634_3;
  wire  T_3634_4;
  wire  T_3634_5;
  wire  T_3634_6;
  wire  T_3634_7;
  wire  T_3634_8;
  wire  T_3634_9;
  wire  T_3634_10;
  wire  T_3634_11;
  wire  T_3634_12;
  wire  T_3634_13;
  wire  T_3634_14;
  wire  T_3634_15;
  wire  T_3634_16;
  wire  T_3639_0;
  wire  T_3639_1;
  wire  T_3639_2;
  wire  T_3639_3;
  wire  T_3639_4;
  wire  T_3639_5;
  wire  T_3639_6;
  wire  T_3639_7;
  wire  T_3639_8;
  wire  T_3639_9;
  wire  T_3639_10;
  wire  T_3639_11;
  wire  T_3639_12;
  wire  T_3639_13;
  wire  T_3639_14;
  wire  T_3639_15;
  wire  T_3639_16;
  wire  T_3644_0;
  wire  T_3644_1;
  wire  T_3644_2;
  wire  T_3644_3;
  wire  T_3644_4;
  wire  T_3644_5;
  wire  T_3644_6;
  wire  T_3644_7;
  wire  T_3644_8;
  wire  T_3644_9;
  wire  T_3644_10;
  wire  T_3644_11;
  wire  T_3644_12;
  wire  T_3644_13;
  wire  T_3644_14;
  wire  T_3644_15;
  wire  T_3644_16;
  wire  T_3806;
  wire  T_3807;
  wire  T_3808;
  wire  T_3809;
  wire [7:0] T_3813;
  wire [7:0] T_3817;
  wire [7:0] T_3821;
  wire [7:0] T_3825;
  wire [15:0] T_3826;
  wire [15:0] T_3827;
  wire [31:0] T_3828;
  wire [31:0] T_3856;
  wire  T_3858;
  wire  T_3911;
  wire [31:0] GEN_7;
  wire  T_3951;
  wire [31:0] GEN_8;
  wire  T_3991;
  wire [31:0] T_4007;
  wire  T_4031;
  wire [31:0] T_4047;
  wire  T_4071;
  wire [31:0] GEN_9;
  wire  T_4111;
  wire [31:0] T_4114;
  wire [31:0] T_4116;
  wire [31:0] T_4117;
  wire [31:0] T_4118;
  wire [31:0] T_4119;
  wire  T_4157;
  wire [31:0] T_4160;
  wire [31:0] T_4162;
  wire [31:0] T_4163;
  wire [31:0] T_4164;
  wire [31:0] T_4165;
  wire  T_4203;
  wire [31:0] T_4219;
  wire  T_4243;
  wire [31:0] GEN_10;
  wire  T_4283;
  wire [31:0] T_4286;
  wire [31:0] T_4288;
  wire [31:0] T_4289;
  wire [31:0] T_4290;
  wire [31:0] T_4291;
  wire  T_4329;
  wire [31:0] GEN_11;
  wire  T_4369;
  wire [31:0] GEN_12;
  wire  T_4409;
  wire [31:0] T_4412;
  wire [31:0] T_4414;
  wire [31:0] T_4415;
  wire [31:0] T_4416;
  wire [31:0] T_4417;
  wire  T_4455;
  wire [31:0] GEN_13;
  wire  T_4495;
  wire [31:0] T_4511;
  wire  T_4535;
  wire [31:0] GEN_14;
  wire  T_4557;
  wire  T_4559;
  wire  T_4561;
  wire  T_4563;
  wire  T_4565;
  wire  T_4567;
  wire  T_4569;
  wire  T_4571;
  wire  T_4573;
  wire  T_4575;
  wire  T_4577;
  wire  T_4579;
  wire  T_4581;
  wire  T_4583;
  wire  T_4585;
  wire  T_4587;
  wire  T_4589;
  wire  T_4591;
  wire  T_4593;
  wire  T_4595;
  wire  T_4597;
  wire  T_4599;
  wire  T_4601;
  wire  T_4603;
  wire  T_4605;
  wire  T_4607;
  wire  T_4609;
  wire  T_4611;
  wire  T_4613;
  wire  T_4615;
  wire  T_4617;
  wire  T_4619;
  wire  T_4621;
  wire  T_4623;
  wire  T_4704_0;
  wire  T_4704_1;
  wire  T_4704_2;
  wire  T_4704_3;
  wire  T_4704_4;
  wire  T_4704_5;
  wire  T_4704_6;
  wire  T_4704_7;
  wire  T_4704_8;
  wire  T_4704_9;
  wire  T_4704_10;
  wire  T_4704_11;
  wire  T_4704_12;
  wire  T_4704_13;
  wire  T_4704_14;
  wire  T_4704_15;
  wire  T_4704_16;
  wire  T_4704_17;
  wire  T_4704_18;
  wire  T_4704_19;
  wire  T_4704_20;
  wire  T_4704_21;
  wire  T_4704_22;
  wire  T_4704_23;
  wire  T_4704_24;
  wire  T_4704_25;
  wire  T_4704_26;
  wire  T_4704_27;
  wire  T_4704_28;
  wire  T_4704_29;
  wire  T_4704_30;
  wire  T_4704_31;
  wire  T_4742;
  wire  T_4746;
  wire  T_4750;
  wire  T_4754;
  wire  T_4758;
  wire  T_4762;
  wire  T_4766;
  wire  T_4770;
  wire  T_4774;
  wire  T_4778;
  wire  T_4782;
  wire  T_4786;
  wire  T_4790;
  wire  T_4794;
  wire  T_4798;
  wire  T_4802;
  wire  T_4806;
  wire  T_4887_0;
  wire  T_4887_1;
  wire  T_4887_2;
  wire  T_4887_3;
  wire  T_4887_4;
  wire  T_4887_5;
  wire  T_4887_6;
  wire  T_4887_7;
  wire  T_4887_8;
  wire  T_4887_9;
  wire  T_4887_10;
  wire  T_4887_11;
  wire  T_4887_12;
  wire  T_4887_13;
  wire  T_4887_14;
  wire  T_4887_15;
  wire  T_4887_16;
  wire  T_4887_17;
  wire  T_4887_18;
  wire  T_4887_19;
  wire  T_4887_20;
  wire  T_4887_21;
  wire  T_4887_22;
  wire  T_4887_23;
  wire  T_4887_24;
  wire  T_4887_25;
  wire  T_4887_26;
  wire  T_4887_27;
  wire  T_4887_28;
  wire  T_4887_29;
  wire  T_4887_30;
  wire  T_4887_31;
  wire  T_4925;
  wire  T_4929;
  wire  T_4933;
  wire  T_4937;
  wire  T_4941;
  wire  T_4945;
  wire  T_4949;
  wire  T_4953;
  wire  T_4957;
  wire  T_4961;
  wire  T_4965;
  wire  T_4969;
  wire  T_4973;
  wire  T_4977;
  wire  T_4981;
  wire  T_4985;
  wire  T_4989;
  wire  T_5070_0;
  wire  T_5070_1;
  wire  T_5070_2;
  wire  T_5070_3;
  wire  T_5070_4;
  wire  T_5070_5;
  wire  T_5070_6;
  wire  T_5070_7;
  wire  T_5070_8;
  wire  T_5070_9;
  wire  T_5070_10;
  wire  T_5070_11;
  wire  T_5070_12;
  wire  T_5070_13;
  wire  T_5070_14;
  wire  T_5070_15;
  wire  T_5070_16;
  wire  T_5070_17;
  wire  T_5070_18;
  wire  T_5070_19;
  wire  T_5070_20;
  wire  T_5070_21;
  wire  T_5070_22;
  wire  T_5070_23;
  wire  T_5070_24;
  wire  T_5070_25;
  wire  T_5070_26;
  wire  T_5070_27;
  wire  T_5070_28;
  wire  T_5070_29;
  wire  T_5070_30;
  wire  T_5070_31;
  wire  T_5108;
  wire  T_5112;
  wire  T_5116;
  wire  T_5120;
  wire  T_5124;
  wire  T_5128;
  wire  T_5132;
  wire  T_5136;
  wire  T_5140;
  wire  T_5144;
  wire  T_5148;
  wire  T_5152;
  wire  T_5156;
  wire  T_5160;
  wire  T_5164;
  wire  T_5168;
  wire  T_5172;
  wire  T_5253_0;
  wire  T_5253_1;
  wire  T_5253_2;
  wire  T_5253_3;
  wire  T_5253_4;
  wire  T_5253_5;
  wire  T_5253_6;
  wire  T_5253_7;
  wire  T_5253_8;
  wire  T_5253_9;
  wire  T_5253_10;
  wire  T_5253_11;
  wire  T_5253_12;
  wire  T_5253_13;
  wire  T_5253_14;
  wire  T_5253_15;
  wire  T_5253_16;
  wire  T_5253_17;
  wire  T_5253_18;
  wire  T_5253_19;
  wire  T_5253_20;
  wire  T_5253_21;
  wire  T_5253_22;
  wire  T_5253_23;
  wire  T_5253_24;
  wire  T_5253_25;
  wire  T_5253_26;
  wire  T_5253_27;
  wire  T_5253_28;
  wire  T_5253_29;
  wire  T_5253_30;
  wire  T_5253_31;
  wire  T_5288;
  wire  T_5289;
  wire  T_5290;
  wire  T_5291;
  wire  T_5292;
  wire [1:0] T_5298;
  wire [1:0] T_5299;
  wire [2:0] T_5300;
  wire [4:0] T_5301;
  wire  GEN_0;
  wire  GEN_15;
  wire  GEN_16;
  wire  GEN_17;
  wire  GEN_18;
  wire  GEN_19;
  wire  GEN_20;
  wire  GEN_21;
  wire  GEN_22;
  wire  GEN_23;
  wire  GEN_24;
  wire  GEN_25;
  wire  GEN_26;
  wire  GEN_27;
  wire  GEN_28;
  wire  GEN_29;
  wire  GEN_30;
  wire  GEN_31;
  wire  GEN_32;
  wire  GEN_33;
  wire  GEN_34;
  wire  GEN_35;
  wire  GEN_36;
  wire  GEN_37;
  wire  GEN_38;
  wire  GEN_39;
  wire  GEN_40;
  wire  GEN_41;
  wire  GEN_42;
  wire  GEN_43;
  wire  GEN_44;
  wire  GEN_45;
  wire  GEN_1;
  wire  GEN_46;
  wire  GEN_47;
  wire  GEN_48;
  wire  GEN_49;
  wire  GEN_50;
  wire  GEN_51;
  wire  GEN_52;
  wire  GEN_53;
  wire  GEN_54;
  wire  GEN_55;
  wire  GEN_56;
  wire  GEN_57;
  wire  GEN_58;
  wire  GEN_59;
  wire  GEN_60;
  wire  GEN_61;
  wire  GEN_62;
  wire  GEN_63;
  wire  GEN_64;
  wire  GEN_65;
  wire  GEN_66;
  wire  GEN_67;
  wire  GEN_68;
  wire  GEN_69;
  wire  GEN_70;
  wire  GEN_71;
  wire  GEN_72;
  wire  GEN_73;
  wire  GEN_74;
  wire  GEN_75;
  wire  GEN_76;
  wire  T_5318;
  wire  GEN_2;
  wire  GEN_77;
  wire  GEN_78;
  wire  GEN_79;
  wire  GEN_80;
  wire  GEN_81;
  wire  GEN_82;
  wire  GEN_83;
  wire  GEN_84;
  wire  GEN_85;
  wire  GEN_86;
  wire  GEN_87;
  wire  GEN_88;
  wire  GEN_89;
  wire  GEN_90;
  wire  GEN_91;
  wire  GEN_92;
  wire  GEN_93;
  wire  GEN_94;
  wire  GEN_95;
  wire  GEN_96;
  wire  GEN_97;
  wire  GEN_98;
  wire  GEN_99;
  wire  GEN_100;
  wire  GEN_101;
  wire  GEN_102;
  wire  GEN_103;
  wire  GEN_104;
  wire  GEN_105;
  wire  GEN_106;
  wire  GEN_107;
  wire  GEN_3;
  wire  GEN_108;
  wire  GEN_109;
  wire  GEN_110;
  wire  GEN_111;
  wire  GEN_112;
  wire  GEN_113;
  wire  GEN_114;
  wire  GEN_115;
  wire  GEN_116;
  wire  GEN_117;
  wire  GEN_118;
  wire  GEN_119;
  wire  GEN_120;
  wire  GEN_121;
  wire  GEN_122;
  wire  GEN_123;
  wire  GEN_124;
  wire  GEN_125;
  wire  GEN_126;
  wire  GEN_127;
  wire  GEN_128;
  wire  GEN_129;
  wire  GEN_130;
  wire  GEN_131;
  wire  GEN_132;
  wire  GEN_133;
  wire  GEN_134;
  wire  GEN_135;
  wire  GEN_136;
  wire  GEN_137;
  wire  GEN_138;
  wire  T_5321;
  wire  T_5322;
  wire  T_5323;
  wire  T_5324;
  wire  T_5325;
  wire [31:0] T_5327;
  wire [1:0] T_5328;
  wire [1:0] T_5329;
  wire [3:0] T_5330;
  wire [1:0] T_5331;
  wire [1:0] T_5332;
  wire [3:0] T_5333;
  wire [7:0] T_5334;
  wire [1:0] T_5335;
  wire [1:0] T_5336;
  wire [3:0] T_5337;
  wire [1:0] T_5338;
  wire [1:0] T_5339;
  wire [3:0] T_5340;
  wire [7:0] T_5341;
  wire [15:0] T_5342;
  wire [1:0] T_5343;
  wire [3:0] T_5345;
  wire [7:0] T_5349;
  wire [15:0] T_5357;
  wire [31:0] T_5358;
  wire [31:0] T_5359;
  wire  T_5394;
  wire  T_5395;
  wire  T_5396;
  wire  T_5397;
  wire  T_5400;
  wire  T_5401;
  wire  T_5403;
  wire  T_5404;
  wire  T_5405;
  wire  T_5407;
  wire  T_5411;
  wire  T_5413;
  wire  T_5416;
  wire  T_5417;
  wire  T_5423;
  wire  T_5427;
  wire  T_5433;
  wire  T_5436;
  wire  T_5437;
  wire  T_5443;
  wire  T_5447;
  wire  T_5453;
  wire  T_5456;
  wire  T_5457;
  wire  T_5463;
  wire  T_5467;
  wire  T_5473;
  wire  T_5476;
  wire  T_5477;
  wire  T_5483;
  wire  T_5487;
  wire  T_5493;
  wire  T_5496;
  wire  T_5497;
  wire  T_5503;
  wire  T_5507;
  wire  T_5513;
  wire  T_5516;
  wire  T_5517;
  wire  T_5523;
  wire  T_5527;
  wire  T_5533;
  wire  T_5536;
  wire  T_5537;
  wire  T_5543;
  wire  T_5547;
  wire  T_5553;
  wire  T_5556;
  wire  T_5557;
  wire  T_5563;
  wire  T_5567;
  wire  T_5573;
  wire  T_5576;
  wire  T_5577;
  wire  T_5583;
  wire  T_5587;
  wire  T_5593;
  wire  T_5596;
  wire  T_5597;
  wire  T_5603;
  wire  T_5607;
  wire  T_5613;
  wire  T_5616;
  wire  T_5617;
  wire  T_5623;
  wire  T_5627;
  wire  T_5633;
  wire  T_5636;
  wire  T_5637;
  wire  T_5643;
  wire  T_5647;
  wire  T_5653;
  wire  T_5656;
  wire  T_5657;
  wire  T_5663;
  wire  T_5667;
  wire  T_5673;
  wire  T_5676;
  wire  T_5677;
  wire  T_5683;
  wire  T_5687;
  wire  T_5693;
  wire  T_5696;
  wire  T_5697;
  wire  T_5703;
  wire  T_5707;
  wire  T_5713;
  wire  T_5716;
  wire  T_5717;
  wire  T_5723;
  wire  T_5727;
  wire  T_5733;
  wire  T_6137_0;
  wire  T_6137_1;
  wire  T_6137_2;
  wire  T_6137_3;
  wire  T_6137_4;
  wire  T_6137_5;
  wire  T_6137_6;
  wire  T_6137_7;
  wire  T_6137_8;
  wire  T_6137_9;
  wire  T_6137_10;
  wire  T_6137_11;
  wire  T_6137_12;
  wire  T_6137_13;
  wire  T_6137_14;
  wire  T_6137_15;
  wire  T_6137_16;
  wire  T_6137_17;
  wire  T_6137_18;
  wire  T_6137_19;
  wire  T_6137_20;
  wire  T_6137_21;
  wire  T_6137_22;
  wire  T_6137_23;
  wire  T_6137_24;
  wire  T_6137_25;
  wire  T_6137_26;
  wire  T_6137_27;
  wire  T_6137_28;
  wire  T_6137_29;
  wire  T_6137_30;
  wire  T_6137_31;
  wire [31:0] T_6208_0;
  wire [31:0] T_6208_1;
  wire [31:0] T_6208_2;
  wire [31:0] T_6208_3;
  wire [31:0] T_6208_4;
  wire [31:0] T_6208_5;
  wire [31:0] T_6208_6;
  wire [31:0] T_6208_7;
  wire [31:0] T_6208_8;
  wire [31:0] T_6208_9;
  wire [31:0] T_6208_10;
  wire [31:0] T_6208_11;
  wire [31:0] T_6208_12;
  wire [31:0] T_6208_13;
  wire [31:0] T_6208_14;
  wire [31:0] T_6208_15;
  wire [31:0] T_6208_16;
  wire [31:0] T_6208_17;
  wire [31:0] T_6208_18;
  wire [31:0] T_6208_19;
  wire [31:0] T_6208_20;
  wire [31:0] T_6208_21;
  wire [31:0] T_6208_22;
  wire [31:0] T_6208_23;
  wire [31:0] T_6208_24;
  wire [31:0] T_6208_25;
  wire [31:0] T_6208_26;
  wire [31:0] T_6208_27;
  wire [31:0] T_6208_28;
  wire [31:0] T_6208_29;
  wire [31:0] T_6208_30;
  wire [31:0] T_6208_31;
  wire  GEN_4;
  wire  GEN_139;
  wire  GEN_140;
  wire  GEN_141;
  wire  GEN_142;
  wire  GEN_143;
  wire  GEN_144;
  wire  GEN_145;
  wire  GEN_146;
  wire  GEN_147;
  wire  GEN_148;
  wire  GEN_149;
  wire  GEN_150;
  wire  GEN_151;
  wire  GEN_152;
  wire  GEN_153;
  wire  GEN_154;
  wire  GEN_155;
  wire  GEN_156;
  wire  GEN_157;
  wire  GEN_158;
  wire  GEN_159;
  wire  GEN_160;
  wire  GEN_161;
  wire  GEN_162;
  wire  GEN_163;
  wire  GEN_164;
  wire  GEN_165;
  wire  GEN_166;
  wire  GEN_167;
  wire  GEN_168;
  wire  GEN_169;
  wire [31:0] GEN_5;
  wire [31:0] GEN_170;
  wire [31:0] GEN_171;
  wire [31:0] GEN_172;
  wire [31:0] GEN_173;
  wire [31:0] GEN_174;
  wire [31:0] GEN_175;
  wire [31:0] GEN_176;
  wire [31:0] GEN_177;
  wire [31:0] GEN_178;
  wire [31:0] GEN_179;
  wire [31:0] GEN_180;
  wire [31:0] GEN_181;
  wire [31:0] GEN_182;
  wire [31:0] GEN_183;
  wire [31:0] GEN_184;
  wire [31:0] GEN_185;
  wire [31:0] GEN_186;
  wire [31:0] GEN_187;
  wire [31:0] GEN_188;
  wire [31:0] GEN_189;
  wire [31:0] GEN_190;
  wire [31:0] GEN_191;
  wire [31:0] GEN_192;
  wire [31:0] GEN_193;
  wire [31:0] GEN_194;
  wire [31:0] GEN_195;
  wire [31:0] GEN_196;
  wire [31:0] GEN_197;
  wire [31:0] GEN_198;
  wire [31:0] GEN_199;
  wire [31:0] GEN_200;
  wire [31:0] T_6245;
  wire [1:0] T_6246;
  wire [4:0] T_6248;
  wire [2:0] T_6249;
  wire [2:0] T_6260_opcode;
  wire [1:0] T_6260_param;
  wire [2:0] T_6260_size;
  wire [4:0] T_6260_source;
  wire  T_6260_sink;
  wire [1:0] T_6260_addr_lo;
  wire [31:0] T_6260_data;
  wire  T_6260_error;
  wire  swPinCtrl_0_oval;
  wire  swPinCtrl_0_oe;
  wire  swPinCtrl_0_ie;
  wire  swPinCtrl_0_pue;
  wire  swPinCtrl_0_ds;
  wire  swPinCtrl_1_oval;
  wire  swPinCtrl_1_oe;
  wire  swPinCtrl_1_ie;
  wire  swPinCtrl_1_pue;
  wire  swPinCtrl_1_ds;
  wire  swPinCtrl_2_oval;
  wire  swPinCtrl_2_oe;
  wire  swPinCtrl_2_ie;
  wire  swPinCtrl_2_pue;
  wire  swPinCtrl_2_ds;
  wire  swPinCtrl_3_oval;
  wire  swPinCtrl_3_oe;
  wire  swPinCtrl_3_ie;
  wire  swPinCtrl_3_pue;
  wire  swPinCtrl_3_ds;
  wire  swPinCtrl_4_oval;
  wire  swPinCtrl_4_oe;
  wire  swPinCtrl_4_ie;
  wire  swPinCtrl_4_pue;
  wire  swPinCtrl_4_ds;
  wire  swPinCtrl_5_oval;
  wire  swPinCtrl_5_oe;
  wire  swPinCtrl_5_ie;
  wire  swPinCtrl_5_pue;
  wire  swPinCtrl_5_ds;
  wire  swPinCtrl_6_oval;
  wire  swPinCtrl_6_oe;
  wire  swPinCtrl_6_ie;
  wire  swPinCtrl_6_pue;
  wire  swPinCtrl_6_ds;
  wire  swPinCtrl_7_oval;
  wire  swPinCtrl_7_oe;
  wire  swPinCtrl_7_ie;
  wire  swPinCtrl_7_pue;
  wire  swPinCtrl_7_ds;
  wire  swPinCtrl_8_oval;
  wire  swPinCtrl_8_oe;
  wire  swPinCtrl_8_ie;
  wire  swPinCtrl_8_pue;
  wire  swPinCtrl_8_ds;
  wire  swPinCtrl_9_oval;
  wire  swPinCtrl_9_oe;
  wire  swPinCtrl_9_ie;
  wire  swPinCtrl_9_pue;
  wire  swPinCtrl_9_ds;
  wire  swPinCtrl_10_oval;
  wire  swPinCtrl_10_oe;
  wire  swPinCtrl_10_ie;
  wire  swPinCtrl_10_pue;
  wire  swPinCtrl_10_ds;
  wire  swPinCtrl_11_oval;
  wire  swPinCtrl_11_oe;
  wire  swPinCtrl_11_ie;
  wire  swPinCtrl_11_pue;
  wire  swPinCtrl_11_ds;
  wire  swPinCtrl_12_oval;
  wire  swPinCtrl_12_oe;
  wire  swPinCtrl_12_ie;
  wire  swPinCtrl_12_pue;
  wire  swPinCtrl_12_ds;
  wire  swPinCtrl_13_oval;
  wire  swPinCtrl_13_oe;
  wire  swPinCtrl_13_ie;
  wire  swPinCtrl_13_pue;
  wire  swPinCtrl_13_ds;
  wire  swPinCtrl_14_oval;
  wire  swPinCtrl_14_oe;
  wire  swPinCtrl_14_ie;
  wire  swPinCtrl_14_pue;
  wire  swPinCtrl_14_ds;
  wire  swPinCtrl_15_oval;
  wire  swPinCtrl_15_oe;
  wire  swPinCtrl_15_ie;
  wire  swPinCtrl_15_pue;
  wire  swPinCtrl_15_ds;
  wire  swPinCtrl_16_oval;
  wire  swPinCtrl_16_oe;
  wire  swPinCtrl_16_ie;
  wire  swPinCtrl_16_pue;
  wire  swPinCtrl_16_ds;
  wire  swPinCtrl_17_oval;
  wire  swPinCtrl_17_oe;
  wire  swPinCtrl_17_ie;
  wire  swPinCtrl_17_pue;
  wire  swPinCtrl_17_ds;
  wire  swPinCtrl_18_oval;
  wire  swPinCtrl_18_oe;
  wire  swPinCtrl_18_ie;
  wire  swPinCtrl_18_pue;
  wire  swPinCtrl_18_ds;
  wire  swPinCtrl_19_oval;
  wire  swPinCtrl_19_oe;
  wire  swPinCtrl_19_ie;
  wire  swPinCtrl_19_pue;
  wire  swPinCtrl_19_ds;
  wire  swPinCtrl_20_oval;
  wire  swPinCtrl_20_oe;
  wire  swPinCtrl_20_ie;
  wire  swPinCtrl_20_pue;
  wire  swPinCtrl_20_ds;
  wire  swPinCtrl_21_oval;
  wire  swPinCtrl_21_oe;
  wire  swPinCtrl_21_ie;
  wire  swPinCtrl_21_pue;
  wire  swPinCtrl_21_ds;
  wire  swPinCtrl_22_oval;
  wire  swPinCtrl_22_oe;
  wire  swPinCtrl_22_ie;
  wire  swPinCtrl_22_pue;
  wire  swPinCtrl_22_ds;
  wire  swPinCtrl_23_oval;
  wire  swPinCtrl_23_oe;
  wire  swPinCtrl_23_ie;
  wire  swPinCtrl_23_pue;
  wire  swPinCtrl_23_ds;
  wire  swPinCtrl_24_oval;
  wire  swPinCtrl_24_oe;
  wire  swPinCtrl_24_ie;
  wire  swPinCtrl_24_pue;
  wire  swPinCtrl_24_ds;
  wire  swPinCtrl_25_oval;
  wire  swPinCtrl_25_oe;
  wire  swPinCtrl_25_ie;
  wire  swPinCtrl_25_pue;
  wire  swPinCtrl_25_ds;
  wire  swPinCtrl_26_oval;
  wire  swPinCtrl_26_oe;
  wire  swPinCtrl_26_ie;
  wire  swPinCtrl_26_pue;
  wire  swPinCtrl_26_ds;
  wire  swPinCtrl_27_oval;
  wire  swPinCtrl_27_oe;
  wire  swPinCtrl_27_ie;
  wire  swPinCtrl_27_pue;
  wire  swPinCtrl_27_ds;
  wire  swPinCtrl_28_oval;
  wire  swPinCtrl_28_oe;
  wire  swPinCtrl_28_ie;
  wire  swPinCtrl_28_pue;
  wire  swPinCtrl_28_ds;
  wire  swPinCtrl_29_oval;
  wire  swPinCtrl_29_oe;
  wire  swPinCtrl_29_ie;
  wire  swPinCtrl_29_pue;
  wire  swPinCtrl_29_ds;
  wire  swPinCtrl_30_oval;
  wire  swPinCtrl_30_oe;
  wire  swPinCtrl_30_ie;
  wire  swPinCtrl_30_pue;
  wire  swPinCtrl_30_ds;
  wire  swPinCtrl_31_oval;
  wire  swPinCtrl_31_oe;
  wire  swPinCtrl_31_ie;
  wire  swPinCtrl_31_pue;
  wire  swPinCtrl_31_ds;
  wire  iof0Ctrl_0_oval;
  wire  iof0Ctrl_0_oe;
  wire  iof0Ctrl_0_ie;
  wire  iof0Ctrl_1_oval;
  wire  iof0Ctrl_1_oe;
  wire  iof0Ctrl_1_ie;
  wire  iof0Ctrl_2_oval;
  wire  iof0Ctrl_2_oe;
  wire  iof0Ctrl_2_ie;
  wire  iof0Ctrl_3_oval;
  wire  iof0Ctrl_3_oe;
  wire  iof0Ctrl_3_ie;
  wire  iof0Ctrl_4_oval;
  wire  iof0Ctrl_4_oe;
  wire  iof0Ctrl_4_ie;
  wire  iof0Ctrl_5_oval;
  wire  iof0Ctrl_5_oe;
  wire  iof0Ctrl_5_ie;
  wire  iof0Ctrl_6_oval;
  wire  iof0Ctrl_6_oe;
  wire  iof0Ctrl_6_ie;
  wire  iof0Ctrl_7_oval;
  wire  iof0Ctrl_7_oe;
  wire  iof0Ctrl_7_ie;
  wire  iof0Ctrl_8_oval;
  wire  iof0Ctrl_8_oe;
  wire  iof0Ctrl_8_ie;
  wire  iof0Ctrl_9_oval;
  wire  iof0Ctrl_9_oe;
  wire  iof0Ctrl_9_ie;
  wire  iof0Ctrl_10_oval;
  wire  iof0Ctrl_10_oe;
  wire  iof0Ctrl_10_ie;
  wire  iof0Ctrl_11_oval;
  wire  iof0Ctrl_11_oe;
  wire  iof0Ctrl_11_ie;
  wire  iof0Ctrl_12_oval;
  wire  iof0Ctrl_12_oe;
  wire  iof0Ctrl_12_ie;
  wire  iof0Ctrl_13_oval;
  wire  iof0Ctrl_13_oe;
  wire  iof0Ctrl_13_ie;
  wire  iof0Ctrl_14_oval;
  wire  iof0Ctrl_14_oe;
  wire  iof0Ctrl_14_ie;
  wire  iof0Ctrl_15_oval;
  wire  iof0Ctrl_15_oe;
  wire  iof0Ctrl_15_ie;
  wire  iof0Ctrl_16_oval;
  wire  iof0Ctrl_16_oe;
  wire  iof0Ctrl_16_ie;
  wire  iof0Ctrl_17_oval;
  wire  iof0Ctrl_17_oe;
  wire  iof0Ctrl_17_ie;
  wire  iof0Ctrl_18_oval;
  wire  iof0Ctrl_18_oe;
  wire  iof0Ctrl_18_ie;
  wire  iof0Ctrl_19_oval;
  wire  iof0Ctrl_19_oe;
  wire  iof0Ctrl_19_ie;
  wire  iof0Ctrl_20_oval;
  wire  iof0Ctrl_20_oe;
  wire  iof0Ctrl_20_ie;
  wire  iof0Ctrl_21_oval;
  wire  iof0Ctrl_21_oe;
  wire  iof0Ctrl_21_ie;
  wire  iof0Ctrl_22_oval;
  wire  iof0Ctrl_22_oe;
  wire  iof0Ctrl_22_ie;
  wire  iof0Ctrl_23_oval;
  wire  iof0Ctrl_23_oe;
  wire  iof0Ctrl_23_ie;
  wire  iof0Ctrl_24_oval;
  wire  iof0Ctrl_24_oe;
  wire  iof0Ctrl_24_ie;
  wire  iof0Ctrl_25_oval;
  wire  iof0Ctrl_25_oe;
  wire  iof0Ctrl_25_ie;
  wire  iof0Ctrl_26_oval;
  wire  iof0Ctrl_26_oe;
  wire  iof0Ctrl_26_ie;
  wire  iof0Ctrl_27_oval;
  wire  iof0Ctrl_27_oe;
  wire  iof0Ctrl_27_ie;
  wire  iof0Ctrl_28_oval;
  wire  iof0Ctrl_28_oe;
  wire  iof0Ctrl_28_ie;
  wire  iof0Ctrl_29_oval;
  wire  iof0Ctrl_29_oe;
  wire  iof0Ctrl_29_ie;
  wire  iof0Ctrl_30_oval;
  wire  iof0Ctrl_30_oe;
  wire  iof0Ctrl_30_ie;
  wire  iof0Ctrl_31_oval;
  wire  iof0Ctrl_31_oe;
  wire  iof0Ctrl_31_ie;
  wire  iof1Ctrl_0_oval;
  wire  iof1Ctrl_0_oe;
  wire  iof1Ctrl_0_ie;
  wire  iof1Ctrl_1_oval;
  wire  iof1Ctrl_1_oe;
  wire  iof1Ctrl_1_ie;
  wire  iof1Ctrl_2_oval;
  wire  iof1Ctrl_2_oe;
  wire  iof1Ctrl_2_ie;
  wire  iof1Ctrl_3_oval;
  wire  iof1Ctrl_3_oe;
  wire  iof1Ctrl_3_ie;
  wire  iof1Ctrl_4_oval;
  wire  iof1Ctrl_4_oe;
  wire  iof1Ctrl_4_ie;
  wire  iof1Ctrl_5_oval;
  wire  iof1Ctrl_5_oe;
  wire  iof1Ctrl_5_ie;
  wire  iof1Ctrl_6_oval;
  wire  iof1Ctrl_6_oe;
  wire  iof1Ctrl_6_ie;
  wire  iof1Ctrl_7_oval;
  wire  iof1Ctrl_7_oe;
  wire  iof1Ctrl_7_ie;
  wire  iof1Ctrl_8_oval;
  wire  iof1Ctrl_8_oe;
  wire  iof1Ctrl_8_ie;
  wire  iof1Ctrl_9_oval;
  wire  iof1Ctrl_9_oe;
  wire  iof1Ctrl_9_ie;
  wire  iof1Ctrl_10_oval;
  wire  iof1Ctrl_10_oe;
  wire  iof1Ctrl_10_ie;
  wire  iof1Ctrl_11_oval;
  wire  iof1Ctrl_11_oe;
  wire  iof1Ctrl_11_ie;
  wire  iof1Ctrl_12_oval;
  wire  iof1Ctrl_12_oe;
  wire  iof1Ctrl_12_ie;
  wire  iof1Ctrl_13_oval;
  wire  iof1Ctrl_13_oe;
  wire  iof1Ctrl_13_ie;
  wire  iof1Ctrl_14_oval;
  wire  iof1Ctrl_14_oe;
  wire  iof1Ctrl_14_ie;
  wire  iof1Ctrl_15_oval;
  wire  iof1Ctrl_15_oe;
  wire  iof1Ctrl_15_ie;
  wire  iof1Ctrl_16_oval;
  wire  iof1Ctrl_16_oe;
  wire  iof1Ctrl_16_ie;
  wire  iof1Ctrl_17_oval;
  wire  iof1Ctrl_17_oe;
  wire  iof1Ctrl_17_ie;
  wire  iof1Ctrl_18_oval;
  wire  iof1Ctrl_18_oe;
  wire  iof1Ctrl_18_ie;
  wire  iof1Ctrl_19_oval;
  wire  iof1Ctrl_19_oe;
  wire  iof1Ctrl_19_ie;
  wire  iof1Ctrl_20_oval;
  wire  iof1Ctrl_20_oe;
  wire  iof1Ctrl_20_ie;
  wire  iof1Ctrl_21_oval;
  wire  iof1Ctrl_21_oe;
  wire  iof1Ctrl_21_ie;
  wire  iof1Ctrl_22_oval;
  wire  iof1Ctrl_22_oe;
  wire  iof1Ctrl_22_ie;
  wire  iof1Ctrl_23_oval;
  wire  iof1Ctrl_23_oe;
  wire  iof1Ctrl_23_ie;
  wire  iof1Ctrl_24_oval;
  wire  iof1Ctrl_24_oe;
  wire  iof1Ctrl_24_ie;
  wire  iof1Ctrl_25_oval;
  wire  iof1Ctrl_25_oe;
  wire  iof1Ctrl_25_ie;
  wire  iof1Ctrl_26_oval;
  wire  iof1Ctrl_26_oe;
  wire  iof1Ctrl_26_ie;
  wire  iof1Ctrl_27_oval;
  wire  iof1Ctrl_27_oe;
  wire  iof1Ctrl_27_ie;
  wire  iof1Ctrl_28_oval;
  wire  iof1Ctrl_28_oe;
  wire  iof1Ctrl_28_ie;
  wire  iof1Ctrl_29_oval;
  wire  iof1Ctrl_29_oe;
  wire  iof1Ctrl_29_ie;
  wire  iof1Ctrl_30_oval;
  wire  iof1Ctrl_30_oe;
  wire  iof1Ctrl_30_ie;
  wire  iof1Ctrl_31_oval;
  wire  iof1Ctrl_31_oe;
  wire  iof1Ctrl_31_ie;
  wire  iofCtrl_0_oval;
  wire  iofCtrl_0_oe;
  wire  iofCtrl_0_ie;
  wire  iofCtrl_1_oval;
  wire  iofCtrl_1_oe;
  wire  iofCtrl_1_ie;
  wire  iofCtrl_2_oval;
  wire  iofCtrl_2_oe;
  wire  iofCtrl_2_ie;
  wire  iofCtrl_3_oval;
  wire  iofCtrl_3_oe;
  wire  iofCtrl_3_ie;
  wire  iofCtrl_4_oval;
  wire  iofCtrl_4_oe;
  wire  iofCtrl_4_ie;
  wire  iofCtrl_5_oval;
  wire  iofCtrl_5_oe;
  wire  iofCtrl_5_ie;
  wire  iofCtrl_6_oval;
  wire  iofCtrl_6_oe;
  wire  iofCtrl_6_ie;
  wire  iofCtrl_7_oval;
  wire  iofCtrl_7_oe;
  wire  iofCtrl_7_ie;
  wire  iofCtrl_8_oval;
  wire  iofCtrl_8_oe;
  wire  iofCtrl_8_ie;
  wire  iofCtrl_9_oval;
  wire  iofCtrl_9_oe;
  wire  iofCtrl_9_ie;
  wire  iofCtrl_10_oval;
  wire  iofCtrl_10_oe;
  wire  iofCtrl_10_ie;
  wire  iofCtrl_11_oval;
  wire  iofCtrl_11_oe;
  wire  iofCtrl_11_ie;
  wire  iofCtrl_12_oval;
  wire  iofCtrl_12_oe;
  wire  iofCtrl_12_ie;
  wire  iofCtrl_13_oval;
  wire  iofCtrl_13_oe;
  wire  iofCtrl_13_ie;
  wire  iofCtrl_14_oval;
  wire  iofCtrl_14_oe;
  wire  iofCtrl_14_ie;
  wire  iofCtrl_15_oval;
  wire  iofCtrl_15_oe;
  wire  iofCtrl_15_ie;
  wire  iofCtrl_16_oval;
  wire  iofCtrl_16_oe;
  wire  iofCtrl_16_ie;
  wire  iofCtrl_17_oval;
  wire  iofCtrl_17_oe;
  wire  iofCtrl_17_ie;
  wire  iofCtrl_18_oval;
  wire  iofCtrl_18_oe;
  wire  iofCtrl_18_ie;
  wire  iofCtrl_19_oval;
  wire  iofCtrl_19_oe;
  wire  iofCtrl_19_ie;
  wire  iofCtrl_20_oval;
  wire  iofCtrl_20_oe;
  wire  iofCtrl_20_ie;
  wire  iofCtrl_21_oval;
  wire  iofCtrl_21_oe;
  wire  iofCtrl_21_ie;
  wire  iofCtrl_22_oval;
  wire  iofCtrl_22_oe;
  wire  iofCtrl_22_ie;
  wire  iofCtrl_23_oval;
  wire  iofCtrl_23_oe;
  wire  iofCtrl_23_ie;
  wire  iofCtrl_24_oval;
  wire  iofCtrl_24_oe;
  wire  iofCtrl_24_ie;
  wire  iofCtrl_25_oval;
  wire  iofCtrl_25_oe;
  wire  iofCtrl_25_ie;
  wire  iofCtrl_26_oval;
  wire  iofCtrl_26_oe;
  wire  iofCtrl_26_ie;
  wire  iofCtrl_27_oval;
  wire  iofCtrl_27_oe;
  wire  iofCtrl_27_ie;
  wire  iofCtrl_28_oval;
  wire  iofCtrl_28_oe;
  wire  iofCtrl_28_ie;
  wire  iofCtrl_29_oval;
  wire  iofCtrl_29_oe;
  wire  iofCtrl_29_ie;
  wire  iofCtrl_30_oval;
  wire  iofCtrl_30_oe;
  wire  iofCtrl_30_ie;
  wire  iofCtrl_31_oval;
  wire  iofCtrl_31_oe;
  wire  iofCtrl_31_ie;
  wire  iofPlusSwPinCtrl_0_oval;
  wire  iofPlusSwPinCtrl_0_oe;
  wire  iofPlusSwPinCtrl_0_ie;
  wire  iofPlusSwPinCtrl_0_pue;
  wire  iofPlusSwPinCtrl_0_ds;
  wire  iofPlusSwPinCtrl_1_oval;
  wire  iofPlusSwPinCtrl_1_oe;
  wire  iofPlusSwPinCtrl_1_ie;
  wire  iofPlusSwPinCtrl_1_pue;
  wire  iofPlusSwPinCtrl_1_ds;
  wire  iofPlusSwPinCtrl_2_oval;
  wire  iofPlusSwPinCtrl_2_oe;
  wire  iofPlusSwPinCtrl_2_ie;
  wire  iofPlusSwPinCtrl_2_pue;
  wire  iofPlusSwPinCtrl_2_ds;
  wire  iofPlusSwPinCtrl_3_oval;
  wire  iofPlusSwPinCtrl_3_oe;
  wire  iofPlusSwPinCtrl_3_ie;
  wire  iofPlusSwPinCtrl_3_pue;
  wire  iofPlusSwPinCtrl_3_ds;
  wire  iofPlusSwPinCtrl_4_oval;
  wire  iofPlusSwPinCtrl_4_oe;
  wire  iofPlusSwPinCtrl_4_ie;
  wire  iofPlusSwPinCtrl_4_pue;
  wire  iofPlusSwPinCtrl_4_ds;
  wire  iofPlusSwPinCtrl_5_oval;
  wire  iofPlusSwPinCtrl_5_oe;
  wire  iofPlusSwPinCtrl_5_ie;
  wire  iofPlusSwPinCtrl_5_pue;
  wire  iofPlusSwPinCtrl_5_ds;
  wire  iofPlusSwPinCtrl_6_oval;
  wire  iofPlusSwPinCtrl_6_oe;
  wire  iofPlusSwPinCtrl_6_ie;
  wire  iofPlusSwPinCtrl_6_pue;
  wire  iofPlusSwPinCtrl_6_ds;
  wire  iofPlusSwPinCtrl_7_oval;
  wire  iofPlusSwPinCtrl_7_oe;
  wire  iofPlusSwPinCtrl_7_ie;
  wire  iofPlusSwPinCtrl_7_pue;
  wire  iofPlusSwPinCtrl_7_ds;
  wire  iofPlusSwPinCtrl_8_oval;
  wire  iofPlusSwPinCtrl_8_oe;
  wire  iofPlusSwPinCtrl_8_ie;
  wire  iofPlusSwPinCtrl_8_pue;
  wire  iofPlusSwPinCtrl_8_ds;
  wire  iofPlusSwPinCtrl_9_oval;
  wire  iofPlusSwPinCtrl_9_oe;
  wire  iofPlusSwPinCtrl_9_ie;
  wire  iofPlusSwPinCtrl_9_pue;
  wire  iofPlusSwPinCtrl_9_ds;
  wire  iofPlusSwPinCtrl_10_oval;
  wire  iofPlusSwPinCtrl_10_oe;
  wire  iofPlusSwPinCtrl_10_ie;
  wire  iofPlusSwPinCtrl_10_pue;
  wire  iofPlusSwPinCtrl_10_ds;
  wire  iofPlusSwPinCtrl_11_oval;
  wire  iofPlusSwPinCtrl_11_oe;
  wire  iofPlusSwPinCtrl_11_ie;
  wire  iofPlusSwPinCtrl_11_pue;
  wire  iofPlusSwPinCtrl_11_ds;
  wire  iofPlusSwPinCtrl_12_oval;
  wire  iofPlusSwPinCtrl_12_oe;
  wire  iofPlusSwPinCtrl_12_ie;
  wire  iofPlusSwPinCtrl_12_pue;
  wire  iofPlusSwPinCtrl_12_ds;
  wire  iofPlusSwPinCtrl_13_oval;
  wire  iofPlusSwPinCtrl_13_oe;
  wire  iofPlusSwPinCtrl_13_ie;
  wire  iofPlusSwPinCtrl_13_pue;
  wire  iofPlusSwPinCtrl_13_ds;
  wire  iofPlusSwPinCtrl_14_oval;
  wire  iofPlusSwPinCtrl_14_oe;
  wire  iofPlusSwPinCtrl_14_ie;
  wire  iofPlusSwPinCtrl_14_pue;
  wire  iofPlusSwPinCtrl_14_ds;
  wire  iofPlusSwPinCtrl_15_oval;
  wire  iofPlusSwPinCtrl_15_oe;
  wire  iofPlusSwPinCtrl_15_ie;
  wire  iofPlusSwPinCtrl_15_pue;
  wire  iofPlusSwPinCtrl_15_ds;
  wire  iofPlusSwPinCtrl_16_oval;
  wire  iofPlusSwPinCtrl_16_oe;
  wire  iofPlusSwPinCtrl_16_ie;
  wire  iofPlusSwPinCtrl_16_pue;
  wire  iofPlusSwPinCtrl_16_ds;
  wire  iofPlusSwPinCtrl_17_oval;
  wire  iofPlusSwPinCtrl_17_oe;
  wire  iofPlusSwPinCtrl_17_ie;
  wire  iofPlusSwPinCtrl_17_pue;
  wire  iofPlusSwPinCtrl_17_ds;
  wire  iofPlusSwPinCtrl_18_oval;
  wire  iofPlusSwPinCtrl_18_oe;
  wire  iofPlusSwPinCtrl_18_ie;
  wire  iofPlusSwPinCtrl_18_pue;
  wire  iofPlusSwPinCtrl_18_ds;
  wire  iofPlusSwPinCtrl_19_oval;
  wire  iofPlusSwPinCtrl_19_oe;
  wire  iofPlusSwPinCtrl_19_ie;
  wire  iofPlusSwPinCtrl_19_pue;
  wire  iofPlusSwPinCtrl_19_ds;
  wire  iofPlusSwPinCtrl_20_oval;
  wire  iofPlusSwPinCtrl_20_oe;
  wire  iofPlusSwPinCtrl_20_ie;
  wire  iofPlusSwPinCtrl_20_pue;
  wire  iofPlusSwPinCtrl_20_ds;
  wire  iofPlusSwPinCtrl_21_oval;
  wire  iofPlusSwPinCtrl_21_oe;
  wire  iofPlusSwPinCtrl_21_ie;
  wire  iofPlusSwPinCtrl_21_pue;
  wire  iofPlusSwPinCtrl_21_ds;
  wire  iofPlusSwPinCtrl_22_oval;
  wire  iofPlusSwPinCtrl_22_oe;
  wire  iofPlusSwPinCtrl_22_ie;
  wire  iofPlusSwPinCtrl_22_pue;
  wire  iofPlusSwPinCtrl_22_ds;
  wire  iofPlusSwPinCtrl_23_oval;
  wire  iofPlusSwPinCtrl_23_oe;
  wire  iofPlusSwPinCtrl_23_ie;
  wire  iofPlusSwPinCtrl_23_pue;
  wire  iofPlusSwPinCtrl_23_ds;
  wire  iofPlusSwPinCtrl_24_oval;
  wire  iofPlusSwPinCtrl_24_oe;
  wire  iofPlusSwPinCtrl_24_ie;
  wire  iofPlusSwPinCtrl_24_pue;
  wire  iofPlusSwPinCtrl_24_ds;
  wire  iofPlusSwPinCtrl_25_oval;
  wire  iofPlusSwPinCtrl_25_oe;
  wire  iofPlusSwPinCtrl_25_ie;
  wire  iofPlusSwPinCtrl_25_pue;
  wire  iofPlusSwPinCtrl_25_ds;
  wire  iofPlusSwPinCtrl_26_oval;
  wire  iofPlusSwPinCtrl_26_oe;
  wire  iofPlusSwPinCtrl_26_ie;
  wire  iofPlusSwPinCtrl_26_pue;
  wire  iofPlusSwPinCtrl_26_ds;
  wire  iofPlusSwPinCtrl_27_oval;
  wire  iofPlusSwPinCtrl_27_oe;
  wire  iofPlusSwPinCtrl_27_ie;
  wire  iofPlusSwPinCtrl_27_pue;
  wire  iofPlusSwPinCtrl_27_ds;
  wire  iofPlusSwPinCtrl_28_oval;
  wire  iofPlusSwPinCtrl_28_oe;
  wire  iofPlusSwPinCtrl_28_ie;
  wire  iofPlusSwPinCtrl_28_pue;
  wire  iofPlusSwPinCtrl_28_ds;
  wire  iofPlusSwPinCtrl_29_oval;
  wire  iofPlusSwPinCtrl_29_oe;
  wire  iofPlusSwPinCtrl_29_ie;
  wire  iofPlusSwPinCtrl_29_pue;
  wire  iofPlusSwPinCtrl_29_ds;
  wire  iofPlusSwPinCtrl_30_oval;
  wire  iofPlusSwPinCtrl_30_oe;
  wire  iofPlusSwPinCtrl_30_ie;
  wire  iofPlusSwPinCtrl_30_pue;
  wire  iofPlusSwPinCtrl_30_ds;
  wire  iofPlusSwPinCtrl_31_oval;
  wire  iofPlusSwPinCtrl_31_oe;
  wire  iofPlusSwPinCtrl_31_ie;
  wire  iofPlusSwPinCtrl_31_pue;
  wire  iofPlusSwPinCtrl_31_ds;
  wire  T_7569;
  wire  T_7570;
  wire  T_7571;
  wire  T_7572;
  wire  T_7573;
  wire  GEN_201;
  wire  GEN_202;
  wire  GEN_203;
  wire  GEN_204;
  wire  GEN_205;
  wire  GEN_206;
  wire  T_7574;
  wire  T_7575_oval;
  wire  T_7575_oe;
  wire  T_7575_ie;
  wire  T_7579;
  wire  T_7580_oval;
  wire  T_7580_oe;
  wire  T_7580_ie;
  wire  T_7580_pue;
  wire  T_7580_ds;
  wire  T_7586;
  wire  T_7587;
  wire  T_7588;
  wire  T_7589;
  wire  T_7590;
  wire  T_7591;
  wire  T_7592;
  wire  T_7593;
  wire  T_7594;
  wire  T_7595;
  wire  T_7596;
  wire  T_7597;
  wire  T_7598;
  wire  T_7599;
  wire  T_7600;
  wire  T_7601;
  wire  T_7602;
  wire  T_7603;
  wire  T_7605;
  wire  T_7606;
  wire  T_7607;
  wire  T_7608;
  wire  T_7609;
  wire  GEN_207;
  wire  GEN_208;
  wire  GEN_209;
  wire  GEN_210;
  wire  GEN_211;
  wire  GEN_212;
  wire  T_7610;
  wire  T_7611_oval;
  wire  T_7611_oe;
  wire  T_7611_ie;
  wire  T_7615;
  wire  T_7616_oval;
  wire  T_7616_oe;
  wire  T_7616_ie;
  wire  T_7616_pue;
  wire  T_7616_ds;
  wire  T_7622;
  wire  T_7623;
  wire  T_7624;
  wire  T_7625;
  wire  T_7626;
  wire  T_7627;
  wire  T_7628;
  wire  T_7629;
  wire  T_7630;
  wire  T_7631;
  wire  T_7632;
  wire  T_7633;
  wire  T_7634;
  wire  T_7635;
  wire  T_7636;
  wire  T_7637;
  wire  T_7638;
  wire  T_7639;
  wire  T_7641;
  wire  T_7642;
  wire  T_7643;
  wire  T_7644;
  wire  T_7645;
  wire  GEN_213;
  wire  GEN_214;
  wire  GEN_215;
  wire  GEN_216;
  wire  GEN_217;
  wire  GEN_218;
  wire  T_7646;
  wire  T_7647_oval;
  wire  T_7647_oe;
  wire  T_7647_ie;
  wire  T_7651;
  wire  T_7652_oval;
  wire  T_7652_oe;
  wire  T_7652_ie;
  wire  T_7652_pue;
  wire  T_7652_ds;
  wire  T_7658;
  wire  T_7659;
  wire  T_7660;
  wire  T_7661;
  wire  T_7662;
  wire  T_7663;
  wire  T_7664;
  wire  T_7665;
  wire  T_7666;
  wire  T_7667;
  wire  T_7668;
  wire  T_7669;
  wire  T_7670;
  wire  T_7671;
  wire  T_7672;
  wire  T_7673;
  wire  T_7674;
  wire  T_7675;
  wire  T_7677;
  wire  T_7678;
  wire  T_7679;
  wire  T_7680;
  wire  T_7681;
  wire  GEN_219;
  wire  GEN_220;
  wire  GEN_221;
  wire  GEN_222;
  wire  GEN_223;
  wire  GEN_224;
  wire  T_7682;
  wire  T_7683_oval;
  wire  T_7683_oe;
  wire  T_7683_ie;
  wire  T_7687;
  wire  T_7688_oval;
  wire  T_7688_oe;
  wire  T_7688_ie;
  wire  T_7688_pue;
  wire  T_7688_ds;
  wire  T_7694;
  wire  T_7695;
  wire  T_7696;
  wire  T_7697;
  wire  T_7698;
  wire  T_7699;
  wire  T_7700;
  wire  T_7701;
  wire  T_7702;
  wire  T_7703;
  wire  T_7704;
  wire  T_7705;
  wire  T_7706;
  wire  T_7707;
  wire  T_7708;
  wire  T_7709;
  wire  T_7710;
  wire  T_7711;
  wire  T_7713;
  wire  T_7714;
  wire  T_7715;
  wire  T_7716;
  wire  T_7717;
  wire  GEN_225;
  wire  GEN_226;
  wire  GEN_227;
  wire  GEN_228;
  wire  GEN_229;
  wire  GEN_230;
  wire  T_7718;
  wire  T_7719_oval;
  wire  T_7719_oe;
  wire  T_7719_ie;
  wire  T_7723;
  wire  T_7724_oval;
  wire  T_7724_oe;
  wire  T_7724_ie;
  wire  T_7724_pue;
  wire  T_7724_ds;
  wire  T_7730;
  wire  T_7731;
  wire  T_7732;
  wire  T_7733;
  wire  T_7734;
  wire  T_7735;
  wire  T_7736;
  wire  T_7737;
  wire  T_7738;
  wire  T_7739;
  wire  T_7740;
  wire  T_7741;
  wire  T_7742;
  wire  T_7743;
  wire  T_7744;
  wire  T_7745;
  wire  T_7746;
  wire  T_7747;
  wire  T_7749;
  wire  T_7750;
  wire  T_7751;
  wire  T_7752;
  wire  T_7753;
  wire  GEN_231;
  wire  GEN_232;
  wire  GEN_233;
  wire  GEN_234;
  wire  GEN_235;
  wire  GEN_236;
  wire  T_7754;
  wire  T_7755_oval;
  wire  T_7755_oe;
  wire  T_7755_ie;
  wire  T_7759;
  wire  T_7760_oval;
  wire  T_7760_oe;
  wire  T_7760_ie;
  wire  T_7760_pue;
  wire  T_7760_ds;
  wire  T_7766;
  wire  T_7767;
  wire  T_7768;
  wire  T_7769;
  wire  T_7770;
  wire  T_7771;
  wire  T_7772;
  wire  T_7773;
  wire  T_7774;
  wire  T_7775;
  wire  T_7776;
  wire  T_7777;
  wire  T_7778;
  wire  T_7779;
  wire  T_7780;
  wire  T_7781;
  wire  T_7782;
  wire  T_7783;
  wire  T_7785;
  wire  T_7786;
  wire  T_7787;
  wire  T_7788;
  wire  T_7789;
  wire  GEN_237;
  wire  GEN_238;
  wire  GEN_239;
  wire  GEN_240;
  wire  GEN_241;
  wire  GEN_242;
  wire  T_7790;
  wire  T_7791_oval;
  wire  T_7791_oe;
  wire  T_7791_ie;
  wire  T_7795;
  wire  T_7796_oval;
  wire  T_7796_oe;
  wire  T_7796_ie;
  wire  T_7796_pue;
  wire  T_7796_ds;
  wire  T_7802;
  wire  T_7803;
  wire  T_7804;
  wire  T_7805;
  wire  T_7806;
  wire  T_7807;
  wire  T_7808;
  wire  T_7809;
  wire  T_7810;
  wire  T_7811;
  wire  T_7812;
  wire  T_7813;
  wire  T_7814;
  wire  T_7815;
  wire  T_7816;
  wire  T_7817;
  wire  T_7818;
  wire  T_7819;
  wire  T_7821;
  wire  T_7822;
  wire  T_7823;
  wire  T_7824;
  wire  T_7825;
  wire  GEN_243;
  wire  GEN_244;
  wire  GEN_245;
  wire  GEN_246;
  wire  GEN_247;
  wire  GEN_248;
  wire  T_7826;
  wire  T_7827_oval;
  wire  T_7827_oe;
  wire  T_7827_ie;
  wire  T_7831;
  wire  T_7832_oval;
  wire  T_7832_oe;
  wire  T_7832_ie;
  wire  T_7832_pue;
  wire  T_7832_ds;
  wire  T_7838;
  wire  T_7839;
  wire  T_7840;
  wire  T_7841;
  wire  T_7842;
  wire  T_7843;
  wire  T_7844;
  wire  T_7845;
  wire  T_7846;
  wire  T_7847;
  wire  T_7848;
  wire  T_7849;
  wire  T_7850;
  wire  T_7851;
  wire  T_7852;
  wire  T_7853;
  wire  T_7854;
  wire  T_7855;
  wire  T_7857;
  wire  T_7858;
  wire  T_7859;
  wire  T_7860;
  wire  T_7861;
  wire  GEN_249;
  wire  GEN_250;
  wire  GEN_251;
  wire  GEN_252;
  wire  GEN_253;
  wire  GEN_254;
  wire  T_7862;
  wire  T_7863_oval;
  wire  T_7863_oe;
  wire  T_7863_ie;
  wire  T_7867;
  wire  T_7868_oval;
  wire  T_7868_oe;
  wire  T_7868_ie;
  wire  T_7868_pue;
  wire  T_7868_ds;
  wire  T_7874;
  wire  T_7875;
  wire  T_7876;
  wire  T_7877;
  wire  T_7878;
  wire  T_7879;
  wire  T_7880;
  wire  T_7881;
  wire  T_7882;
  wire  T_7883;
  wire  T_7884;
  wire  T_7885;
  wire  T_7886;
  wire  T_7887;
  wire  T_7888;
  wire  T_7889;
  wire  T_7890;
  wire  T_7891;
  wire  T_7893;
  wire  T_7894;
  wire  T_7895;
  wire  T_7896;
  wire  T_7897;
  wire  GEN_255;
  wire  GEN_256;
  wire  GEN_257;
  wire  GEN_258;
  wire  GEN_259;
  wire  GEN_260;
  wire  T_7898;
  wire  T_7899_oval;
  wire  T_7899_oe;
  wire  T_7899_ie;
  wire  T_7903;
  wire  T_7904_oval;
  wire  T_7904_oe;
  wire  T_7904_ie;
  wire  T_7904_pue;
  wire  T_7904_ds;
  wire  T_7910;
  wire  T_7911;
  wire  T_7912;
  wire  T_7913;
  wire  T_7914;
  wire  T_7915;
  wire  T_7916;
  wire  T_7917;
  wire  T_7918;
  wire  T_7919;
  wire  T_7920;
  wire  T_7921;
  wire  T_7922;
  wire  T_7923;
  wire  T_7924;
  wire  T_7925;
  wire  T_7926;
  wire  T_7927;
  wire  T_7929;
  wire  T_7930;
  wire  T_7931;
  wire  T_7932;
  wire  T_7933;
  wire  GEN_261;
  wire  GEN_262;
  wire  GEN_263;
  wire  GEN_264;
  wire  GEN_265;
  wire  GEN_266;
  wire  T_7934;
  wire  T_7935_oval;
  wire  T_7935_oe;
  wire  T_7935_ie;
  wire  T_7939;
  wire  T_7940_oval;
  wire  T_7940_oe;
  wire  T_7940_ie;
  wire  T_7940_pue;
  wire  T_7940_ds;
  wire  T_7946;
  wire  T_7947;
  wire  T_7948;
  wire  T_7949;
  wire  T_7950;
  wire  T_7951;
  wire  T_7952;
  wire  T_7953;
  wire  T_7954;
  wire  T_7955;
  wire  T_7956;
  wire  T_7957;
  wire  T_7958;
  wire  T_7959;
  wire  T_7960;
  wire  T_7961;
  wire  T_7962;
  wire  T_7963;
  wire  T_7965;
  wire  T_7966;
  wire  T_7967;
  wire  T_7968;
  wire  T_7969;
  wire  GEN_267;
  wire  GEN_268;
  wire  GEN_269;
  wire  GEN_270;
  wire  GEN_271;
  wire  GEN_272;
  wire  T_7970;
  wire  T_7971_oval;
  wire  T_7971_oe;
  wire  T_7971_ie;
  wire  T_7975;
  wire  T_7976_oval;
  wire  T_7976_oe;
  wire  T_7976_ie;
  wire  T_7976_pue;
  wire  T_7976_ds;
  wire  T_7982;
  wire  T_7983;
  wire  T_7984;
  wire  T_7985;
  wire  T_7986;
  wire  T_7987;
  wire  T_7988;
  wire  T_7989;
  wire  T_7990;
  wire  T_7991;
  wire  T_7992;
  wire  T_7993;
  wire  T_7994;
  wire  T_7995;
  wire  T_7996;
  wire  T_7997;
  wire  T_7998;
  wire  T_7999;
  wire  T_8001;
  wire  T_8002;
  wire  T_8003;
  wire  T_8004;
  wire  T_8005;
  wire  GEN_273;
  wire  GEN_274;
  wire  GEN_275;
  wire  GEN_276;
  wire  GEN_277;
  wire  GEN_278;
  wire  T_8006;
  wire  T_8007_oval;
  wire  T_8007_oe;
  wire  T_8007_ie;
  wire  T_8011;
  wire  T_8012_oval;
  wire  T_8012_oe;
  wire  T_8012_ie;
  wire  T_8012_pue;
  wire  T_8012_ds;
  wire  T_8018;
  wire  T_8019;
  wire  T_8020;
  wire  T_8021;
  wire  T_8022;
  wire  T_8023;
  wire  T_8024;
  wire  T_8025;
  wire  T_8026;
  wire  T_8027;
  wire  T_8028;
  wire  T_8029;
  wire  T_8030;
  wire  T_8031;
  wire  T_8032;
  wire  T_8033;
  wire  T_8034;
  wire  T_8035;
  wire  T_8037;
  wire  T_8038;
  wire  T_8039;
  wire  T_8040;
  wire  T_8041;
  wire  GEN_279;
  wire  GEN_280;
  wire  GEN_281;
  wire  GEN_282;
  wire  GEN_283;
  wire  GEN_284;
  wire  T_8042;
  wire  T_8043_oval;
  wire  T_8043_oe;
  wire  T_8043_ie;
  wire  T_8047;
  wire  T_8048_oval;
  wire  T_8048_oe;
  wire  T_8048_ie;
  wire  T_8048_pue;
  wire  T_8048_ds;
  wire  T_8054;
  wire  T_8055;
  wire  T_8056;
  wire  T_8057;
  wire  T_8058;
  wire  T_8059;
  wire  T_8060;
  wire  T_8061;
  wire  T_8062;
  wire  T_8063;
  wire  T_8064;
  wire  T_8065;
  wire  T_8066;
  wire  T_8067;
  wire  T_8068;
  wire  T_8069;
  wire  T_8070;
  wire  T_8071;
  wire  T_8073;
  wire  T_8074;
  wire  T_8075;
  wire  T_8076;
  wire  T_8077;
  wire  GEN_285;
  wire  GEN_286;
  wire  GEN_287;
  wire  GEN_288;
  wire  GEN_289;
  wire  GEN_290;
  wire  T_8078;
  wire  T_8079_oval;
  wire  T_8079_oe;
  wire  T_8079_ie;
  wire  T_8083;
  wire  T_8084_oval;
  wire  T_8084_oe;
  wire  T_8084_ie;
  wire  T_8084_pue;
  wire  T_8084_ds;
  wire  T_8090;
  wire  T_8091;
  wire  T_8092;
  wire  T_8093;
  wire  T_8094;
  wire  T_8095;
  wire  T_8096;
  wire  T_8097;
  wire  T_8098;
  wire  T_8099;
  wire  T_8100;
  wire  T_8101;
  wire  T_8102;
  wire  T_8103;
  wire  T_8104;
  wire  T_8105;
  wire  T_8106;
  wire  T_8107;
  wire  T_8109;
  wire  T_8110;
  wire  T_8111;
  wire  T_8112;
  wire  T_8113;
  wire  GEN_291;
  wire  GEN_292;
  wire  GEN_293;
  wire  GEN_294;
  wire  GEN_295;
  wire  GEN_296;
  wire  T_8114;
  wire  T_8115_oval;
  wire  T_8115_oe;
  wire  T_8115_ie;
  wire  T_8119;
  wire  T_8120_oval;
  wire  T_8120_oe;
  wire  T_8120_ie;
  wire  T_8120_pue;
  wire  T_8120_ds;
  wire  T_8126;
  wire  T_8127;
  wire  T_8128;
  wire  T_8129;
  wire  T_8130;
  wire  T_8131;
  wire  T_8132;
  wire  T_8133;
  wire  T_8134;
  wire  T_8135;
  wire  T_8136;
  wire  T_8137;
  wire  T_8138;
  wire  T_8139;
  wire  T_8140;
  wire  T_8141;
  wire  T_8142;
  wire  T_8143;
  wire  T_8145;
  wire  T_8146;
  wire  T_8147;
  wire  T_8148;
  wire  T_8149;
  wire  GEN_297;
  wire  GEN_298;
  wire  GEN_299;
  wire  GEN_300;
  wire  GEN_301;
  wire  GEN_302;
  wire  T_8150;
  wire  T_8151_oval;
  wire  T_8151_oe;
  wire  T_8151_ie;
  wire  T_8155;
  wire  T_8156_oval;
  wire  T_8156_oe;
  wire  T_8156_ie;
  wire  T_8156_pue;
  wire  T_8156_ds;
  wire  T_8162;
  wire  T_8163;
  wire  T_8164;
  wire  T_8165;
  wire  T_8166;
  wire  T_8167;
  wire  T_8168;
  wire  T_8169;
  wire  T_8170;
  wire  T_8171;
  wire  T_8172;
  wire  T_8173;
  wire  T_8174;
  wire  T_8175;
  wire  T_8176;
  wire  T_8177;
  wire  T_8178;
  wire  T_8179;
  wire  T_8181;
  wire  T_8182;
  wire  T_8183;
  wire  T_8184;
  wire  T_8185;
  wire  GEN_303;
  wire  GEN_304;
  wire  GEN_305;
  wire  GEN_306;
  wire  GEN_307;
  wire  GEN_308;
  wire  T_8186;
  wire  T_8187_oval;
  wire  T_8187_oe;
  wire  T_8187_ie;
  wire  T_8191;
  wire  T_8192_oval;
  wire  T_8192_oe;
  wire  T_8192_ie;
  wire  T_8192_pue;
  wire  T_8192_ds;
  wire  T_8198;
  wire  T_8199;
  wire  T_8200;
  wire  T_8201;
  wire  T_8202;
  wire  T_8203;
  wire  T_8204;
  wire  T_8205;
  wire  T_8206;
  wire  T_8207;
  wire  T_8208;
  wire  T_8209;
  wire  T_8210;
  wire  T_8211;
  wire  T_8212;
  wire  T_8213;
  wire  T_8214;
  wire  T_8215;
  wire  T_8217;
  wire  T_8218;
  wire  T_8219;
  wire  T_8220;
  wire  T_8221;
  wire  GEN_309;
  wire  GEN_310;
  wire  GEN_311;
  wire  GEN_312;
  wire  GEN_313;
  wire  GEN_314;
  wire  T_8222;
  wire  T_8223_oval;
  wire  T_8223_oe;
  wire  T_8223_ie;
  wire  T_8227;
  wire  T_8228_oval;
  wire  T_8228_oe;
  wire  T_8228_ie;
  wire  T_8228_pue;
  wire  T_8228_ds;
  wire  T_8234;
  wire  T_8235;
  wire  T_8236;
  wire  T_8237;
  wire  T_8238;
  wire  T_8239;
  wire  T_8240;
  wire  T_8241;
  wire  T_8242;
  wire  T_8243;
  wire  T_8244;
  wire  T_8245;
  wire  T_8246;
  wire  T_8247;
  wire  T_8248;
  wire  T_8249;
  wire  T_8250;
  wire  T_8251;
  wire  T_8253;
  wire  T_8254;
  wire  T_8255;
  wire  T_8256;
  wire  T_8257;
  wire  GEN_315;
  wire  GEN_316;
  wire  GEN_317;
  wire  GEN_318;
  wire  GEN_319;
  wire  GEN_320;
  wire  T_8258;
  wire  T_8259_oval;
  wire  T_8259_oe;
  wire  T_8259_ie;
  wire  T_8263;
  wire  T_8264_oval;
  wire  T_8264_oe;
  wire  T_8264_ie;
  wire  T_8264_pue;
  wire  T_8264_ds;
  wire  T_8270;
  wire  T_8271;
  wire  T_8272;
  wire  T_8273;
  wire  T_8274;
  wire  T_8275;
  wire  T_8276;
  wire  T_8277;
  wire  T_8278;
  wire  T_8279;
  wire  T_8280;
  wire  T_8281;
  wire  T_8282;
  wire  T_8283;
  wire  T_8284;
  wire  T_8285;
  wire  T_8286;
  wire  T_8287;
  wire  T_8289;
  wire  T_8290;
  wire  T_8291;
  wire  T_8292;
  wire  T_8293;
  wire  GEN_321;
  wire  GEN_322;
  wire  GEN_323;
  wire  GEN_324;
  wire  GEN_325;
  wire  GEN_326;
  wire  T_8294;
  wire  T_8295_oval;
  wire  T_8295_oe;
  wire  T_8295_ie;
  wire  T_8299;
  wire  T_8300_oval;
  wire  T_8300_oe;
  wire  T_8300_ie;
  wire  T_8300_pue;
  wire  T_8300_ds;
  wire  T_8306;
  wire  T_8307;
  wire  T_8308;
  wire  T_8309;
  wire  T_8310;
  wire  T_8311;
  wire  T_8312;
  wire  T_8313;
  wire  T_8314;
  wire  T_8315;
  wire  T_8316;
  wire  T_8317;
  wire  T_8318;
  wire  T_8319;
  wire  T_8320;
  wire  T_8321;
  wire  T_8322;
  wire  T_8323;
  wire  T_8325;
  wire  T_8326;
  wire  T_8327;
  wire  T_8328;
  wire  T_8329;
  wire  GEN_327;
  wire  GEN_328;
  wire  GEN_329;
  wire  GEN_330;
  wire  GEN_331;
  wire  GEN_332;
  wire  T_8330;
  wire  T_8331_oval;
  wire  T_8331_oe;
  wire  T_8331_ie;
  wire  T_8335;
  wire  T_8336_oval;
  wire  T_8336_oe;
  wire  T_8336_ie;
  wire  T_8336_pue;
  wire  T_8336_ds;
  wire  T_8342;
  wire  T_8343;
  wire  T_8344;
  wire  T_8345;
  wire  T_8346;
  wire  T_8347;
  wire  T_8348;
  wire  T_8349;
  wire  T_8350;
  wire  T_8351;
  wire  T_8352;
  wire  T_8353;
  wire  T_8354;
  wire  T_8355;
  wire  T_8356;
  wire  T_8357;
  wire  T_8358;
  wire  T_8359;
  wire  T_8361;
  wire  T_8362;
  wire  T_8363;
  wire  T_8364;
  wire  T_8365;
  wire  GEN_333;
  wire  GEN_334;
  wire  GEN_335;
  wire  GEN_336;
  wire  GEN_337;
  wire  GEN_338;
  wire  T_8366;
  wire  T_8367_oval;
  wire  T_8367_oe;
  wire  T_8367_ie;
  wire  T_8371;
  wire  T_8372_oval;
  wire  T_8372_oe;
  wire  T_8372_ie;
  wire  T_8372_pue;
  wire  T_8372_ds;
  wire  T_8378;
  wire  T_8379;
  wire  T_8380;
  wire  T_8381;
  wire  T_8382;
  wire  T_8383;
  wire  T_8384;
  wire  T_8385;
  wire  T_8386;
  wire  T_8387;
  wire  T_8388;
  wire  T_8389;
  wire  T_8390;
  wire  T_8391;
  wire  T_8392;
  wire  T_8393;
  wire  T_8394;
  wire  T_8395;
  wire  T_8397;
  wire  T_8398;
  wire  T_8399;
  wire  T_8400;
  wire  T_8401;
  wire  GEN_339;
  wire  GEN_340;
  wire  GEN_341;
  wire  GEN_342;
  wire  GEN_343;
  wire  GEN_344;
  wire  T_8402;
  wire  T_8403_oval;
  wire  T_8403_oe;
  wire  T_8403_ie;
  wire  T_8407;
  wire  T_8408_oval;
  wire  T_8408_oe;
  wire  T_8408_ie;
  wire  T_8408_pue;
  wire  T_8408_ds;
  wire  T_8414;
  wire  T_8415;
  wire  T_8416;
  wire  T_8417;
  wire  T_8418;
  wire  T_8419;
  wire  T_8420;
  wire  T_8421;
  wire  T_8422;
  wire  T_8423;
  wire  T_8424;
  wire  T_8425;
  wire  T_8426;
  wire  T_8427;
  wire  T_8428;
  wire  T_8429;
  wire  T_8430;
  wire  T_8431;
  wire  T_8433;
  wire  T_8434;
  wire  T_8435;
  wire  T_8436;
  wire  T_8437;
  wire  GEN_345;
  wire  GEN_346;
  wire  GEN_347;
  wire  GEN_348;
  wire  GEN_349;
  wire  GEN_350;
  wire  T_8438;
  wire  T_8439_oval;
  wire  T_8439_oe;
  wire  T_8439_ie;
  wire  T_8443;
  wire  T_8444_oval;
  wire  T_8444_oe;
  wire  T_8444_ie;
  wire  T_8444_pue;
  wire  T_8444_ds;
  wire  T_8450;
  wire  T_8451;
  wire  T_8452;
  wire  T_8453;
  wire  T_8454;
  wire  T_8455;
  wire  T_8456;
  wire  T_8457;
  wire  T_8458;
  wire  T_8459;
  wire  T_8460;
  wire  T_8461;
  wire  T_8462;
  wire  T_8463;
  wire  T_8464;
  wire  T_8465;
  wire  T_8466;
  wire  T_8467;
  wire  T_8469;
  wire  T_8470;
  wire  T_8471;
  wire  T_8472;
  wire  T_8473;
  wire  GEN_351;
  wire  GEN_352;
  wire  GEN_353;
  wire  GEN_354;
  wire  GEN_355;
  wire  GEN_356;
  wire  T_8474;
  wire  T_8475_oval;
  wire  T_8475_oe;
  wire  T_8475_ie;
  wire  T_8479;
  wire  T_8480_oval;
  wire  T_8480_oe;
  wire  T_8480_ie;
  wire  T_8480_pue;
  wire  T_8480_ds;
  wire  T_8486;
  wire  T_8487;
  wire  T_8488;
  wire  T_8489;
  wire  T_8490;
  wire  T_8491;
  wire  T_8492;
  wire  T_8493;
  wire  T_8494;
  wire  T_8495;
  wire  T_8496;
  wire  T_8497;
  wire  T_8498;
  wire  T_8499;
  wire  T_8500;
  wire  T_8501;
  wire  T_8502;
  wire  T_8503;
  wire  T_8505;
  wire  T_8506;
  wire  T_8507;
  wire  T_8508;
  wire  T_8509;
  wire  GEN_357;
  wire  GEN_358;
  wire  GEN_359;
  wire  GEN_360;
  wire  GEN_361;
  wire  GEN_362;
  wire  T_8510;
  wire  T_8511_oval;
  wire  T_8511_oe;
  wire  T_8511_ie;
  wire  T_8515;
  wire  T_8516_oval;
  wire  T_8516_oe;
  wire  T_8516_ie;
  wire  T_8516_pue;
  wire  T_8516_ds;
  wire  T_8522;
  wire  T_8523;
  wire  T_8524;
  wire  T_8525;
  wire  T_8526;
  wire  T_8527;
  wire  T_8528;
  wire  T_8529;
  wire  T_8530;
  wire  T_8531;
  wire  T_8532;
  wire  T_8533;
  wire  T_8534;
  wire  T_8535;
  wire  T_8536;
  wire  T_8537;
  wire  T_8538;
  wire  T_8539;
  wire  T_8541;
  wire  T_8542;
  wire  T_8543;
  wire  T_8544;
  wire  T_8545;
  wire  GEN_363;
  wire  GEN_364;
  wire  GEN_365;
  wire  GEN_366;
  wire  GEN_367;
  wire  GEN_368;
  wire  T_8546;
  wire  T_8547_oval;
  wire  T_8547_oe;
  wire  T_8547_ie;
  wire  T_8551;
  wire  T_8552_oval;
  wire  T_8552_oe;
  wire  T_8552_ie;
  wire  T_8552_pue;
  wire  T_8552_ds;
  wire  T_8558;
  wire  T_8559;
  wire  T_8560;
  wire  T_8561;
  wire  T_8562;
  wire  T_8563;
  wire  T_8564;
  wire  T_8565;
  wire  T_8566;
  wire  T_8567;
  wire  T_8568;
  wire  T_8569;
  wire  T_8570;
  wire  T_8571;
  wire  T_8572;
  wire  T_8573;
  wire  T_8574;
  wire  T_8575;
  wire  T_8577;
  wire  T_8578;
  wire  T_8579;
  wire  T_8580;
  wire  T_8581;
  wire  GEN_369;
  wire  GEN_370;
  wire  GEN_371;
  wire  GEN_372;
  wire  GEN_373;
  wire  GEN_374;
  wire  T_8582;
  wire  T_8583_oval;
  wire  T_8583_oe;
  wire  T_8583_ie;
  wire  T_8587;
  wire  T_8588_oval;
  wire  T_8588_oe;
  wire  T_8588_ie;
  wire  T_8588_pue;
  wire  T_8588_ds;
  wire  T_8594;
  wire  T_8595;
  wire  T_8596;
  wire  T_8597;
  wire  T_8598;
  wire  T_8599;
  wire  T_8600;
  wire  T_8601;
  wire  T_8602;
  wire  T_8603;
  wire  T_8604;
  wire  T_8605;
  wire  T_8606;
  wire  T_8607;
  wire  T_8608;
  wire  T_8609;
  wire  T_8610;
  wire  T_8611;
  wire  T_8613;
  wire  T_8614;
  wire  T_8615;
  wire  T_8616;
  wire  T_8617;
  wire  GEN_375;
  wire  GEN_376;
  wire  GEN_377;
  wire  GEN_378;
  wire  GEN_379;
  wire  GEN_380;
  wire  T_8618;
  wire  T_8619_oval;
  wire  T_8619_oe;
  wire  T_8619_ie;
  wire  T_8623;
  wire  T_8624_oval;
  wire  T_8624_oe;
  wire  T_8624_ie;
  wire  T_8624_pue;
  wire  T_8624_ds;
  wire  T_8630;
  wire  T_8631;
  wire  T_8632;
  wire  T_8633;
  wire  T_8634;
  wire  T_8635;
  wire  T_8636;
  wire  T_8637;
  wire  T_8638;
  wire  T_8639;
  wire  T_8640;
  wire  T_8641;
  wire  T_8642;
  wire  T_8643;
  wire  T_8644;
  wire  T_8645;
  wire  T_8646;
  wire  T_8647;
  wire  T_8649;
  wire  T_8650;
  wire  T_8651;
  wire  T_8652;
  wire  T_8653;
  wire  GEN_381;
  wire  GEN_382;
  wire  GEN_383;
  wire  GEN_384;
  wire  GEN_385;
  wire  GEN_386;
  wire  T_8654;
  wire  T_8655_oval;
  wire  T_8655_oe;
  wire  T_8655_ie;
  wire  T_8659;
  wire  T_8660_oval;
  wire  T_8660_oe;
  wire  T_8660_ie;
  wire  T_8660_pue;
  wire  T_8660_ds;
  wire  T_8666;
  wire  T_8667;
  wire  T_8668;
  wire  T_8669;
  wire  T_8670;
  wire  T_8671;
  wire  T_8672;
  wire  T_8673;
  wire  T_8674;
  wire  T_8675;
  wire  T_8676;
  wire  T_8677;
  wire  T_8678;
  wire  T_8679;
  wire  T_8680;
  wire  T_8681;
  wire  T_8682;
  wire  T_8683;
  wire  T_8685;
  wire  T_8686;
  wire  T_8687;
  wire  T_8688;
  wire  T_8689;
  wire  GEN_387;
  wire  GEN_388;
  wire  GEN_389;
  wire  GEN_390;
  wire  GEN_391;
  wire  GEN_392;
  wire  T_8690;
  wire  T_8691_oval;
  wire  T_8691_oe;
  wire  T_8691_ie;
  wire  T_8695;
  wire  T_8696_oval;
  wire  T_8696_oe;
  wire  T_8696_ie;
  wire  T_8696_pue;
  wire  T_8696_ds;
  wire  T_8702;
  wire  T_8703;
  wire  T_8704;
  wire  T_8705;
  wire  T_8706;
  wire  T_8707;
  wire  T_8708;
  wire  T_8709;
  wire  T_8710;
  wire  T_8711;
  wire  T_8712;
  wire  T_8713;
  wire  T_8714;
  wire  T_8715;
  wire  T_8716;
  wire  T_8717;
  wire  T_8718;
  wire  T_8719;
  wire [2:0] GEN_6 = 3'b0;
  wire [1:0] GEN_393 = 2'b0;
  wire [2:0] GEN_394 = 3'b0;
  wire [4:0] GEN_395 = 5'b0;
  wire [28:0] GEN_396 = 29'b0;
  wire [3:0] GEN_397 = 4'b0;
  wire [31:0] GEN_398 = 32'b0;
  sirv_AsyncResetRegVec_67 u_oeReg (
    .clock(oeReg_clock),
    .reset(oeReg_reset),
    .io_d(oeReg_io_d),
    .io_q(oeReg_io_q),
    .io_en(oeReg_io_en)
  );
  sirv_AsyncResetRegVec_67 u_pueReg (
    .clock(pueReg_clock),
    .reset(pueReg_reset),
    .io_d(pueReg_io_d),
    .io_q(pueReg_io_q),
    .io_en(pueReg_io_en)
  );
  sirv_AsyncResetRegVec_67 u_ieReg (
    .clock(ieReg_clock),
    .reset(ieReg_reset),
    .io_d(ieReg_io_d),
    .io_q(ieReg_io_q),
    .io_en(ieReg_io_en)
  );
  sirv_AsyncResetRegVec_67 u_iofEnReg (
    .clock(iofEnReg_clock),
    .reset(iofEnReg_reset),
    .io_d(iofEnReg_io_d),
    .io_q(iofEnReg_io_q),
    .io_en(iofEnReg_io_en)
  );
  assign io_interrupts_0_0 = T_7602;
  assign io_interrupts_0_1 = T_7638;
  assign io_interrupts_0_2 = T_7674;
  assign io_interrupts_0_3 = T_7710;
  assign io_interrupts_0_4 = T_7746;
  assign io_interrupts_0_5 = T_7782;
  assign io_interrupts_0_6 = T_7818;
  assign io_interrupts_0_7 = T_7854;
  assign io_interrupts_0_8 = T_7890;
  assign io_interrupts_0_9 = T_7926;
  assign io_interrupts_0_10 = T_7962;
  assign io_interrupts_0_11 = T_7998;
  assign io_interrupts_0_12 = T_8034;
  assign io_interrupts_0_13 = T_8070;
  assign io_interrupts_0_14 = T_8106;
  assign io_interrupts_0_15 = T_8142;
  assign io_interrupts_0_16 = T_8178;
  assign io_interrupts_0_17 = T_8214;
  assign io_interrupts_0_18 = T_8250;
  assign io_interrupts_0_19 = T_8286;
  assign io_interrupts_0_20 = T_8322;
  assign io_interrupts_0_21 = T_8358;
  assign io_interrupts_0_22 = T_8394;
  assign io_interrupts_0_23 = T_8430;
  assign io_interrupts_0_24 = T_8466;
  assign io_interrupts_0_25 = T_8502;
  assign io_interrupts_0_26 = T_8538;
  assign io_interrupts_0_27 = T_8574;
  assign io_interrupts_0_28 = T_8610;
  assign io_interrupts_0_29 = T_8646;
  assign io_interrupts_0_30 = T_8682;
  assign io_interrupts_0_31 = T_8718;
  assign io_in_0_a_ready = T_3295_ready;
  assign io_in_0_b_valid = 1'h0;
  assign io_in_0_b_bits_opcode = GEN_6;
  assign io_in_0_b_bits_param = GEN_393;
  assign io_in_0_b_bits_size = GEN_394;
  assign io_in_0_b_bits_source = GEN_395;
  assign io_in_0_b_bits_address = GEN_396;
  assign io_in_0_b_bits_mask = GEN_397;
  assign io_in_0_b_bits_data = GEN_398;
  assign io_in_0_c_ready = 1'h1;
  assign io_in_0_d_valid = T_3334_valid;
  assign io_in_0_d_bits_opcode = {{2'd0}, T_3334_bits_read};
  assign io_in_0_d_bits_param = T_6260_param;
  assign io_in_0_d_bits_size = T_6260_size;
  assign io_in_0_d_bits_source = T_6260_source;
  assign io_in_0_d_bits_sink = T_6260_sink;
  assign io_in_0_d_bits_addr_lo = T_6260_addr_lo;
  assign io_in_0_d_bits_data = T_3334_bits_data;
  assign io_in_0_d_bits_error = T_6260_error;
  assign io_in_0_e_ready = 1'h1;
  assign io_port_pins_0_o_oval = T_7587;
  assign io_port_pins_0_o_oe = T_7580_oe;
  assign io_port_pins_0_o_ie = T_7580_ie;
  assign io_port_pins_0_o_pue = T_7580_pue;
  assign io_port_pins_0_o_ds = T_7580_ds;
  assign io_port_pins_1_o_oval = T_7623;
  assign io_port_pins_1_o_oe = T_7616_oe;
  assign io_port_pins_1_o_ie = T_7616_ie;
  assign io_port_pins_1_o_pue = T_7616_pue;
  assign io_port_pins_1_o_ds = T_7616_ds;
  assign io_port_pins_2_o_oval = T_7659;
  assign io_port_pins_2_o_oe = T_7652_oe;
  assign io_port_pins_2_o_ie = T_7652_ie;
  assign io_port_pins_2_o_pue = T_7652_pue;
  assign io_port_pins_2_o_ds = T_7652_ds;
  assign io_port_pins_3_o_oval = T_7695;
  assign io_port_pins_3_o_oe = T_7688_oe;
  assign io_port_pins_3_o_ie = T_7688_ie;
  assign io_port_pins_3_o_pue = T_7688_pue;
  assign io_port_pins_3_o_ds = T_7688_ds;
  assign io_port_pins_4_o_oval = T_7731;
  assign io_port_pins_4_o_oe = T_7724_oe;
  assign io_port_pins_4_o_ie = T_7724_ie;
  assign io_port_pins_4_o_pue = T_7724_pue;
  assign io_port_pins_4_o_ds = T_7724_ds;
  assign io_port_pins_5_o_oval = T_7767;
  assign io_port_pins_5_o_oe = T_7760_oe;
  assign io_port_pins_5_o_ie = T_7760_ie;
  assign io_port_pins_5_o_pue = T_7760_pue;
  assign io_port_pins_5_o_ds = T_7760_ds;
  assign io_port_pins_6_o_oval = T_7803;
  assign io_port_pins_6_o_oe = T_7796_oe;
  assign io_port_pins_6_o_ie = T_7796_ie;
  assign io_port_pins_6_o_pue = T_7796_pue;
  assign io_port_pins_6_o_ds = T_7796_ds;
  assign io_port_pins_7_o_oval = T_7839;
  assign io_port_pins_7_o_oe = T_7832_oe;
  assign io_port_pins_7_o_ie = T_7832_ie;
  assign io_port_pins_7_o_pue = T_7832_pue;
  assign io_port_pins_7_o_ds = T_7832_ds;
  assign io_port_pins_8_o_oval = T_7875;
  assign io_port_pins_8_o_oe = T_7868_oe;
  assign io_port_pins_8_o_ie = T_7868_ie;
  assign io_port_pins_8_o_pue = T_7868_pue;
  assign io_port_pins_8_o_ds = T_7868_ds;
  assign io_port_pins_9_o_oval = T_7911;
  assign io_port_pins_9_o_oe = T_7904_oe;
  assign io_port_pins_9_o_ie = T_7904_ie;
  assign io_port_pins_9_o_pue = T_7904_pue;
  assign io_port_pins_9_o_ds = T_7904_ds;
  assign io_port_pins_10_o_oval = T_7947;
  assign io_port_pins_10_o_oe = T_7940_oe;
  assign io_port_pins_10_o_ie = T_7940_ie;
  assign io_port_pins_10_o_pue = T_7940_pue;
  assign io_port_pins_10_o_ds = T_7940_ds;
  assign io_port_pins_11_o_oval = T_7983;
  assign io_port_pins_11_o_oe = T_7976_oe;
  assign io_port_pins_11_o_ie = T_7976_ie;
  assign io_port_pins_11_o_pue = T_7976_pue;
  assign io_port_pins_11_o_ds = T_7976_ds;
  assign io_port_pins_12_o_oval = T_8019;
  assign io_port_pins_12_o_oe = T_8012_oe;
  assign io_port_pins_12_o_ie = T_8012_ie;
  assign io_port_pins_12_o_pue = T_8012_pue;
  assign io_port_pins_12_o_ds = T_8012_ds;
  assign io_port_pins_13_o_oval = T_8055;
  assign io_port_pins_13_o_oe = T_8048_oe;
  assign io_port_pins_13_o_ie = T_8048_ie;
  assign io_port_pins_13_o_pue = T_8048_pue;
  assign io_port_pins_13_o_ds = T_8048_ds;
  assign io_port_pins_14_o_oval = T_8091;
  assign io_port_pins_14_o_oe = T_8084_oe;
  assign io_port_pins_14_o_ie = T_8084_ie;
  assign io_port_pins_14_o_pue = T_8084_pue;
  assign io_port_pins_14_o_ds = T_8084_ds;
  assign io_port_pins_15_o_oval = T_8127;
  assign io_port_pins_15_o_oe = T_8120_oe;
  assign io_port_pins_15_o_ie = T_8120_ie;
  assign io_port_pins_15_o_pue = T_8120_pue;
  assign io_port_pins_15_o_ds = T_8120_ds;
  assign io_port_pins_16_o_oval = T_8163;
  assign io_port_pins_16_o_oe = T_8156_oe;
  assign io_port_pins_16_o_ie = T_8156_ie;
  assign io_port_pins_16_o_pue = T_8156_pue;
  assign io_port_pins_16_o_ds = T_8156_ds;
  assign io_port_pins_17_o_oval = T_8199;
  assign io_port_pins_17_o_oe = T_8192_oe;
  assign io_port_pins_17_o_ie = T_8192_ie;
  assign io_port_pins_17_o_pue = T_8192_pue;
  assign io_port_pins_17_o_ds = T_8192_ds;
  assign io_port_pins_18_o_oval = T_8235;
  assign io_port_pins_18_o_oe = T_8228_oe;
  assign io_port_pins_18_o_ie = T_8228_ie;
  assign io_port_pins_18_o_pue = T_8228_pue;
  assign io_port_pins_18_o_ds = T_8228_ds;
  assign io_port_pins_19_o_oval = T_8271;
  assign io_port_pins_19_o_oe = T_8264_oe;
  assign io_port_pins_19_o_ie = T_8264_ie;
  assign io_port_pins_19_o_pue = T_8264_pue;
  assign io_port_pins_19_o_ds = T_8264_ds;
  assign io_port_pins_20_o_oval = T_8307;
  assign io_port_pins_20_o_oe = T_8300_oe;
  assign io_port_pins_20_o_ie = T_8300_ie;
  assign io_port_pins_20_o_pue = T_8300_pue;
  assign io_port_pins_20_o_ds = T_8300_ds;
  assign io_port_pins_21_o_oval = T_8343;
  assign io_port_pins_21_o_oe = T_8336_oe;
  assign io_port_pins_21_o_ie = T_8336_ie;
  assign io_port_pins_21_o_pue = T_8336_pue;
  assign io_port_pins_21_o_ds = T_8336_ds;
  assign io_port_pins_22_o_oval = T_8379;
  assign io_port_pins_22_o_oe = T_8372_oe;
  assign io_port_pins_22_o_ie = T_8372_ie;
  assign io_port_pins_22_o_pue = T_8372_pue;
  assign io_port_pins_22_o_ds = T_8372_ds;
  assign io_port_pins_23_o_oval = T_8415;
  assign io_port_pins_23_o_oe = T_8408_oe;
  assign io_port_pins_23_o_ie = T_8408_ie;
  assign io_port_pins_23_o_pue = T_8408_pue;
  assign io_port_pins_23_o_ds = T_8408_ds;
  assign io_port_pins_24_o_oval = T_8451;
  assign io_port_pins_24_o_oe = T_8444_oe;
  assign io_port_pins_24_o_ie = T_8444_ie;
  assign io_port_pins_24_o_pue = T_8444_pue;
  assign io_port_pins_24_o_ds = T_8444_ds;
  assign io_port_pins_25_o_oval = T_8487;
  assign io_port_pins_25_o_oe = T_8480_oe;
  assign io_port_pins_25_o_ie = T_8480_ie;
  assign io_port_pins_25_o_pue = T_8480_pue;
  assign io_port_pins_25_o_ds = T_8480_ds;
  assign io_port_pins_26_o_oval = T_8523;
  assign io_port_pins_26_o_oe = T_8516_oe;
  assign io_port_pins_26_o_ie = T_8516_ie;
  assign io_port_pins_26_o_pue = T_8516_pue;
  assign io_port_pins_26_o_ds = T_8516_ds;
  assign io_port_pins_27_o_oval = T_8559;
  assign io_port_pins_27_o_oe = T_8552_oe;
  assign io_port_pins_27_o_ie = T_8552_ie;
  assign io_port_pins_27_o_pue = T_8552_pue;
  assign io_port_pins_27_o_ds = T_8552_ds;
  assign io_port_pins_28_o_oval = T_8595;
  assign io_port_pins_28_o_oe = T_8588_oe;
  assign io_port_pins_28_o_ie = T_8588_ie;
  assign io_port_pins_28_o_pue = T_8588_pue;
  assign io_port_pins_28_o_ds = T_8588_ds;
  assign io_port_pins_29_o_oval = T_8631;
  assign io_port_pins_29_o_oe = T_8624_oe;
  assign io_port_pins_29_o_ie = T_8624_ie;
  assign io_port_pins_29_o_pue = T_8624_pue;
  assign io_port_pins_29_o_ds = T_8624_ds;
  assign io_port_pins_30_o_oval = T_8667;
  assign io_port_pins_30_o_oe = T_8660_oe;
  assign io_port_pins_30_o_ie = T_8660_ie;
  assign io_port_pins_30_o_pue = T_8660_pue;
  assign io_port_pins_30_o_ds = T_8660_ds;
  assign io_port_pins_31_o_oval = T_8703;
  assign io_port_pins_31_o_oe = T_8696_oe;
  assign io_port_pins_31_o_ie = T_8696_ie;
  assign io_port_pins_31_o_pue = T_8696_pue;
  assign io_port_pins_31_o_ds = T_8696_ds;
  assign io_port_iof_0_0_i_ival = T_7603;
  assign io_port_iof_0_1_i_ival = T_7639;
  assign io_port_iof_0_2_i_ival = T_7675;
  assign io_port_iof_0_3_i_ival = T_7711;
  assign io_port_iof_0_4_i_ival = T_7747;
  assign io_port_iof_0_5_i_ival = T_7783;
  assign io_port_iof_0_6_i_ival = T_7819;
  assign io_port_iof_0_7_i_ival = T_7855;
  assign io_port_iof_0_8_i_ival = T_7891;
  assign io_port_iof_0_9_i_ival = T_7927;
  assign io_port_iof_0_10_i_ival = T_7963;
  assign io_port_iof_0_11_i_ival = T_7999;
  assign io_port_iof_0_12_i_ival = T_8035;
  assign io_port_iof_0_13_i_ival = T_8071;
  assign io_port_iof_0_14_i_ival = T_8107;
  assign io_port_iof_0_15_i_ival = T_8143;
  assign io_port_iof_0_16_i_ival = T_8179;
  assign io_port_iof_0_17_i_ival = T_8215;
  assign io_port_iof_0_18_i_ival = T_8251;
  assign io_port_iof_0_19_i_ival = T_8287;
  assign io_port_iof_0_20_i_ival = T_8323;
  assign io_port_iof_0_21_i_ival = T_8359;
  assign io_port_iof_0_22_i_ival = T_8395;
  assign io_port_iof_0_23_i_ival = T_8431;
  assign io_port_iof_0_24_i_ival = T_8467;
  assign io_port_iof_0_25_i_ival = T_8503;
  assign io_port_iof_0_26_i_ival = T_8539;
  assign io_port_iof_0_27_i_ival = T_8575;
  assign io_port_iof_0_28_i_ival = T_8611;
  assign io_port_iof_0_29_i_ival = T_8647;
  assign io_port_iof_0_30_i_ival = T_8683;
  assign io_port_iof_0_31_i_ival = T_8719;
  assign io_port_iof_1_0_i_ival = T_7603;
  assign io_port_iof_1_1_i_ival = T_7639;
  assign io_port_iof_1_2_i_ival = T_7675;
  assign io_port_iof_1_3_i_ival = T_7711;
  assign io_port_iof_1_4_i_ival = T_7747;
  assign io_port_iof_1_5_i_ival = T_7783;
  assign io_port_iof_1_6_i_ival = T_7819;
  assign io_port_iof_1_7_i_ival = T_7855;
  assign io_port_iof_1_8_i_ival = T_7891;
  assign io_port_iof_1_9_i_ival = T_7927;
  assign io_port_iof_1_10_i_ival = T_7963;
  assign io_port_iof_1_11_i_ival = T_7999;
  assign io_port_iof_1_12_i_ival = T_8035;
  assign io_port_iof_1_13_i_ival = T_8071;
  assign io_port_iof_1_14_i_ival = T_8107;
  assign io_port_iof_1_15_i_ival = T_8143;
  assign io_port_iof_1_16_i_ival = T_8179;
  assign io_port_iof_1_17_i_ival = T_8215;
  assign io_port_iof_1_18_i_ival = T_8251;
  assign io_port_iof_1_19_i_ival = T_8287;
  assign io_port_iof_1_20_i_ival = T_8323;
  assign io_port_iof_1_21_i_ival = T_8359;
  assign io_port_iof_1_22_i_ival = T_8395;
  assign io_port_iof_1_23_i_ival = T_8431;
  assign io_port_iof_1_24_i_ival = T_8467;
  assign io_port_iof_1_25_i_ival = T_8503;
  assign io_port_iof_1_26_i_ival = T_8539;
  assign io_port_iof_1_27_i_ival = T_8575;
  assign io_port_iof_1_28_i_ival = T_8611;
  assign io_port_iof_1_29_i_ival = T_8647;
  assign io_port_iof_1_30_i_ival = T_8683;
  assign io_port_iof_1_31_i_ival = T_8719;
  assign oeReg_clock = clock;
  assign oeReg_reset = reset;
  assign oeReg_io_d = T_3370_bits_data;
  assign oeReg_io_en = T_4203;
  assign pueReg_clock = clock;
  assign pueReg_reset = reset;
  assign pueReg_io_d = T_3370_bits_data;
  assign pueReg_io_en = T_4495;
  assign ieReg_clock = clock;
  assign ieReg_reset = reset;
  assign ieReg_io_d = T_3370_bits_data;
  assign ieReg_io_en = T_4031;
  assign inVal = T_3253;
  assign T_3188_0 = io_port_pins_0_i_ival;
  assign T_3188_1 = io_port_pins_1_i_ival;
  assign T_3188_2 = io_port_pins_2_i_ival;
  assign T_3188_3 = io_port_pins_3_i_ival;
  assign T_3188_4 = io_port_pins_4_i_ival;
  assign T_3188_5 = io_port_pins_5_i_ival;
  assign T_3188_6 = io_port_pins_6_i_ival;
  assign T_3188_7 = io_port_pins_7_i_ival;
  assign T_3188_8 = io_port_pins_8_i_ival;
  assign T_3188_9 = io_port_pins_9_i_ival;
  assign T_3188_10 = io_port_pins_10_i_ival;
  assign T_3188_11 = io_port_pins_11_i_ival;
  assign T_3188_12 = io_port_pins_12_i_ival;
  assign T_3188_13 = io_port_pins_13_i_ival;
  assign T_3188_14 = io_port_pins_14_i_ival;
  assign T_3188_15 = io_port_pins_15_i_ival;
  assign T_3188_16 = io_port_pins_16_i_ival;
  assign T_3188_17 = io_port_pins_17_i_ival;
  assign T_3188_18 = io_port_pins_18_i_ival;
  assign T_3188_19 = io_port_pins_19_i_ival;
  assign T_3188_20 = io_port_pins_20_i_ival;
  assign T_3188_21 = io_port_pins_21_i_ival;
  assign T_3188_22 = io_port_pins_22_i_ival;
  assign T_3188_23 = io_port_pins_23_i_ival;
  assign T_3188_24 = io_port_pins_24_i_ival;
  assign T_3188_25 = io_port_pins_25_i_ival;
  assign T_3188_26 = io_port_pins_26_i_ival;
  assign T_3188_27 = io_port_pins_27_i_ival;
  assign T_3188_28 = io_port_pins_28_i_ival;
  assign T_3188_29 = io_port_pins_29_i_ival;
  assign T_3188_30 = io_port_pins_30_i_ival;
  assign T_3188_31 = io_port_pins_31_i_ival;
  assign T_3223 = {T_3188_1,T_3188_0};
  assign T_3224 = {T_3188_3,T_3188_2};
  assign T_3225 = {T_3224,T_3223};
  assign T_3226 = {T_3188_5,T_3188_4};
  assign T_3227 = {T_3188_7,T_3188_6};
  assign T_3228 = {T_3227,T_3226};
  assign T_3229 = {T_3228,T_3225};
  assign T_3230 = {T_3188_9,T_3188_8};
  assign T_3231 = {T_3188_11,T_3188_10};
  assign T_3232 = {T_3231,T_3230};
  assign T_3233 = {T_3188_13,T_3188_12};
  assign T_3234 = {T_3188_15,T_3188_14};
  assign T_3235 = {T_3234,T_3233};
  assign T_3236 = {T_3235,T_3232};
  assign T_3237 = {T_3236,T_3229};
  assign T_3238 = {T_3188_17,T_3188_16};
  assign T_3239 = {T_3188_19,T_3188_18};
  assign T_3240 = {T_3239,T_3238};
  assign T_3241 = {T_3188_21,T_3188_20};
  assign T_3242 = {T_3188_23,T_3188_22};
  assign T_3243 = {T_3242,T_3241};
  assign T_3244 = {T_3243,T_3240};
  assign T_3245 = {T_3188_25,T_3188_24};
  assign T_3246 = {T_3188_27,T_3188_26};
  assign T_3247 = {T_3246,T_3245};
  assign T_3248 = {T_3188_29,T_3188_28};
  assign T_3249 = {T_3188_31,T_3188_30};
  assign T_3250 = {T_3249,T_3248};
  assign T_3251 = {T_3250,T_3247};
  assign T_3252 = {T_3251,T_3244};
  assign T_3253 = {T_3252,T_3237};
  assign iofEnReg_clock = clock;
  assign iofEnReg_reset = reset;
  assign iofEnReg_io_d = T_3370_bits_data;
  assign iofEnReg_io_en = T_3991;
  assign T_3269 = ~ valueReg;
  assign rise = T_3269 & inSyncReg;
  assign T_3270 = ~ inSyncReg;
  assign fall = valueReg & T_3270;
  assign T_3295_ready = T_5322;
  assign T_3295_valid = io_in_0_a_valid;
  assign T_3295_bits_read = T_3312;
  assign T_3295_bits_index = T_3313[9:0];
  assign T_3295_bits_data = io_in_0_a_bits_data;
  assign T_3295_bits_mask = io_in_0_a_bits_mask;
  assign T_3295_bits_extra = T_3316;
  assign T_3312 = io_in_0_a_bits_opcode == 3'h4;
  assign T_3313 = io_in_0_a_bits_address[28:2];
  assign T_3314 = io_in_0_a_bits_address[1:0];
  assign T_3315 = {T_3314,io_in_0_a_bits_source};
  assign T_3316 = {T_3315,io_in_0_a_bits_size};
  assign T_3334_ready = io_in_0_d_ready;
  assign T_3334_valid = T_5325;
  assign T_3334_bits_read = T_3370_bits_read;
  assign T_3334_bits_data = T_6245;
  assign T_3334_bits_extra = T_3370_bits_extra;
  assign T_3370_ready = T_5324;
  assign T_3370_valid = T_5323;
  assign T_3370_bits_read = T_3295_bits_read;
  assign T_3370_bits_index = T_3295_bits_index;
  assign T_3370_bits_data = T_3295_bits_data;
  assign T_3370_bits_mask = T_3295_bits_mask;
  assign T_3370_bits_extra = T_3295_bits_extra;
  assign T_3455 = T_3370_bits_index & 10'h3e0;
  assign T_3457 = T_3455 == 10'h0;
  assign T_3463 = T_3370_bits_index ^ 10'h5;
  assign T_3464 = T_3463 & 10'h3e0;
  assign T_3466 = T_3464 == 10'h0;
  assign T_3472 = T_3370_bits_index ^ 10'ha;
  assign T_3473 = T_3472 & 10'h3e0;
  assign T_3475 = T_3473 == 10'h0;
  assign T_3481 = T_3370_bits_index ^ 10'he;
  assign T_3482 = T_3481 & 10'h3e0;
  assign T_3484 = T_3482 == 10'h0;
  assign T_3490 = T_3370_bits_index ^ 10'h1;
  assign T_3491 = T_3490 & 10'h3e0;
  assign T_3493 = T_3491 == 10'h0;
  assign T_3499 = T_3370_bits_index ^ 10'h6;
  assign T_3500 = T_3499 & 10'h3e0;
  assign T_3502 = T_3500 == 10'h0;
  assign T_3508 = T_3370_bits_index ^ 10'h9;
  assign T_3509 = T_3508 & 10'h3e0;
  assign T_3511 = T_3509 == 10'h0;
  assign T_3517 = T_3370_bits_index ^ 10'hd;
  assign T_3518 = T_3517 & 10'h3e0;
  assign T_3520 = T_3518 == 10'h0;
  assign T_3526 = T_3370_bits_index ^ 10'h2;
  assign T_3527 = T_3526 & 10'h3e0;
  assign T_3529 = T_3527 == 10'h0;
  assign T_3535 = T_3370_bits_index ^ 10'hc;
  assign T_3536 = T_3535 & 10'h3e0;
  assign T_3538 = T_3536 == 10'h0;
  assign T_3544 = T_3370_bits_index ^ 10'h7;
  assign T_3545 = T_3544 & 10'h3e0;
  assign T_3547 = T_3545 == 10'h0;
  assign T_3553 = T_3370_bits_index ^ 10'h3;
  assign T_3554 = T_3553 & 10'h3e0;
  assign T_3556 = T_3554 == 10'h0;
  assign T_3562 = T_3370_bits_index ^ 10'h10;
  assign T_3563 = T_3562 & 10'h3e0;
  assign T_3565 = T_3563 == 10'h0;
  assign T_3571 = T_3370_bits_index ^ 10'hb;
  assign T_3572 = T_3571 & 10'h3e0;
  assign T_3574 = T_3572 == 10'h0;
  assign T_3580 = T_3370_bits_index ^ 10'h8;
  assign T_3581 = T_3580 & 10'h3e0;
  assign T_3583 = T_3581 == 10'h0;
  assign T_3589 = T_3370_bits_index ^ 10'h4;
  assign T_3590 = T_3589 & 10'h3e0;
  assign T_3592 = T_3590 == 10'h0;
  assign T_3598 = T_3370_bits_index ^ 10'hf;
  assign T_3599 = T_3598 & 10'h3e0;
  assign T_3601 = T_3599 == 10'h0;
  assign T_3609_0 = T_5397;
  assign T_3609_1 = T_5497;
  assign T_3609_2 = T_5597;
  assign T_3609_3 = T_5677;
  assign T_3609_4 = T_5417;
  assign T_3609_5 = T_5517;
  assign T_3609_6 = T_5577;
  assign T_3609_7 = T_5657;
  assign T_3609_8 = T_5437;
  assign T_3609_9 = T_5637;
  assign T_3609_10 = T_5537;
  assign T_3609_11 = T_5457;
  assign T_3609_12 = T_5717;
  assign T_3609_13 = T_5617;
  assign T_3609_14 = T_5557;
  assign T_3609_15 = T_5477;
  assign T_3609_16 = T_5697;
  assign T_3614_0 = T_5403;
  assign T_3614_1 = T_5503;
  assign T_3614_2 = T_5603;
  assign T_3614_3 = T_5683;
  assign T_3614_4 = T_5423;
  assign T_3614_5 = T_5523;
  assign T_3614_6 = T_5583;
  assign T_3614_7 = T_5663;
  assign T_3614_8 = T_5443;
  assign T_3614_9 = T_5643;
  assign T_3614_10 = T_5543;
  assign T_3614_11 = T_5463;
  assign T_3614_12 = T_5723;
  assign T_3614_13 = T_5623;
  assign T_3614_14 = T_5563;
  assign T_3614_15 = T_5483;
  assign T_3614_16 = T_5703;
  assign T_3619_0 = 1'h1;
  assign T_3619_1 = 1'h1;
  assign T_3619_2 = 1'h1;
  assign T_3619_3 = 1'h1;
  assign T_3619_4 = 1'h1;
  assign T_3619_5 = 1'h1;
  assign T_3619_6 = 1'h1;
  assign T_3619_7 = 1'h1;
  assign T_3619_8 = 1'h1;
  assign T_3619_9 = 1'h1;
  assign T_3619_10 = 1'h1;
  assign T_3619_11 = 1'h1;
  assign T_3619_12 = 1'h1;
  assign T_3619_13 = 1'h1;
  assign T_3619_14 = 1'h1;
  assign T_3619_15 = 1'h1;
  assign T_3619_16 = 1'h1;
  assign T_3624_0 = 1'h1;
  assign T_3624_1 = 1'h1;
  assign T_3624_2 = 1'h1;
  assign T_3624_3 = 1'h1;
  assign T_3624_4 = 1'h1;
  assign T_3624_5 = 1'h1;
  assign T_3624_6 = 1'h1;
  assign T_3624_7 = 1'h1;
  assign T_3624_8 = 1'h1;
  assign T_3624_9 = 1'h1;
  assign T_3624_10 = 1'h1;
  assign T_3624_11 = 1'h1;
  assign T_3624_12 = 1'h1;
  assign T_3624_13 = 1'h1;
  assign T_3624_14 = 1'h1;
  assign T_3624_15 = 1'h1;
  assign T_3624_16 = 1'h1;
  assign T_3629_0 = 1'h1;
  assign T_3629_1 = 1'h1;
  assign T_3629_2 = 1'h1;
  assign T_3629_3 = 1'h1;
  assign T_3629_4 = 1'h1;
  assign T_3629_5 = 1'h1;
  assign T_3629_6 = 1'h1;
  assign T_3629_7 = 1'h1;
  assign T_3629_8 = 1'h1;
  assign T_3629_9 = 1'h1;
  assign T_3629_10 = 1'h1;
  assign T_3629_11 = 1'h1;
  assign T_3629_12 = 1'h1;
  assign T_3629_13 = 1'h1;
  assign T_3629_14 = 1'h1;
  assign T_3629_15 = 1'h1;
  assign T_3629_16 = 1'h1;
  assign T_3634_0 = 1'h1;
  assign T_3634_1 = 1'h1;
  assign T_3634_2 = 1'h1;
  assign T_3634_3 = 1'h1;
  assign T_3634_4 = 1'h1;
  assign T_3634_5 = 1'h1;
  assign T_3634_6 = 1'h1;
  assign T_3634_7 = 1'h1;
  assign T_3634_8 = 1'h1;
  assign T_3634_9 = 1'h1;
  assign T_3634_10 = 1'h1;
  assign T_3634_11 = 1'h1;
  assign T_3634_12 = 1'h1;
  assign T_3634_13 = 1'h1;
  assign T_3634_14 = 1'h1;
  assign T_3634_15 = 1'h1;
  assign T_3634_16 = 1'h1;
  assign T_3639_0 = T_5407;
  assign T_3639_1 = T_5507;
  assign T_3639_2 = T_5607;
  assign T_3639_3 = T_5687;
  assign T_3639_4 = T_5427;
  assign T_3639_5 = T_5527;
  assign T_3639_6 = T_5587;
  assign T_3639_7 = T_5667;
  assign T_3639_8 = T_5447;
  assign T_3639_9 = T_5647;
  assign T_3639_10 = T_5547;
  assign T_3639_11 = T_5467;
  assign T_3639_12 = T_5727;
  assign T_3639_13 = T_5627;
  assign T_3639_14 = T_5567;
  assign T_3639_15 = T_5487;
  assign T_3639_16 = T_5707;
  assign T_3644_0 = T_5413;
  assign T_3644_1 = T_5513;
  assign T_3644_2 = T_5613;
  assign T_3644_3 = T_5693;
  assign T_3644_4 = T_5433;
  assign T_3644_5 = T_5533;
  assign T_3644_6 = T_5593;
  assign T_3644_7 = T_5673;
  assign T_3644_8 = T_5453;
  assign T_3644_9 = T_5653;
  assign T_3644_10 = T_5553;
  assign T_3644_11 = T_5473;
  assign T_3644_12 = T_5733;
  assign T_3644_13 = T_5633;
  assign T_3644_14 = T_5573;
  assign T_3644_15 = T_5493;
  assign T_3644_16 = T_5713;
  assign T_3806 = T_3370_bits_mask[0];
  assign T_3807 = T_3370_bits_mask[1];
  assign T_3808 = T_3370_bits_mask[2];
  assign T_3809 = T_3370_bits_mask[3];
  assign T_3813 = T_3806 ? 8'hff : 8'h0;
  assign T_3817 = T_3807 ? 8'hff : 8'h0;
  assign T_3821 = T_3808 ? 8'hff : 8'h0;
  assign T_3825 = T_3809 ? 8'hff : 8'h0;
  assign T_3826 = {T_3817,T_3813};
  assign T_3827 = {T_3825,T_3821};
  assign T_3828 = {T_3827,T_3826};
  assign T_3856 = ~ T_3828;
  assign T_3858 = T_3856 == 32'h0;
  assign T_3911 = T_3644_1 & T_3858;
  assign GEN_7 = T_3911 ? T_3370_bits_data : dsReg;
  assign T_3951 = T_3644_2 & T_3858;
  assign GEN_8 = T_3951 ? T_3370_bits_data : highIeReg;
  assign T_3991 = T_3644_3 & T_3858;
  assign T_4007 = iofEnReg_io_q;
  assign T_4031 = T_3644_4 & T_3858;
  assign T_4047 = ieReg_io_q;
  assign T_4071 = T_3644_5 & T_3858;
  assign GEN_9 = T_4071 ? T_3370_bits_data : riseIeReg;
  assign T_4111 = T_3644_6 & T_3858;
  assign T_4114 = ~ fallIpReg;
  assign T_4116 = T_4111 ? T_3370_bits_data : 32'h0;
  assign T_4117 = T_4114 | T_4116;
  assign T_4118 = ~ T_4117;
  assign T_4119 = T_4118 | fall;
  assign T_4157 = T_3644_7 & T_3858;
  assign T_4160 = ~ lowIpReg;
  assign T_4162 = T_4157 ? T_3370_bits_data : 32'h0;
  assign T_4163 = T_4160 | T_4162;
  assign T_4164 = ~ T_4163;
  assign T_4165 = T_4164 | T_3269;
  assign T_4203 = T_3644_8 & T_3858;
  assign T_4219 = oeReg_io_q;
  assign T_4243 = T_3644_9 & T_3858;
  assign GEN_10 = T_4243 ? T_3370_bits_data : lowIeReg;
  assign T_4283 = T_3644_10 & T_3858;
  assign T_4286 = ~ riseIpReg;
  assign T_4288 = T_4283 ? T_3370_bits_data : 32'h0;
  assign T_4289 = T_4286 | T_4288;
  assign T_4290 = ~ T_4289;
  assign T_4291 = T_4290 | rise;
  assign T_4329 = T_3644_11 & T_3858;
  assign GEN_11 = T_4329 ? T_3370_bits_data : portReg;
  assign T_4369 = T_3644_12 & T_3858;
  assign GEN_12 = T_4369 ? T_3370_bits_data : xorReg;
  assign T_4409 = T_3644_13 & T_3858;
  assign T_4412 = ~ highIpReg;
  assign T_4414 = T_4409 ? T_3370_bits_data : 32'h0;
  assign T_4415 = T_4412 | T_4414;
  assign T_4416 = ~ T_4415;
  assign T_4417 = T_4416 | valueReg;
  assign T_4455 = T_3644_14 & T_3858;
  assign GEN_13 = T_4455 ? T_3370_bits_data : fallIeReg;
  assign T_4495 = T_3644_15 & T_3858;
  assign T_4511 = pueReg_io_q;
  assign T_4535 = T_3644_16 & T_3858;
  assign GEN_14 = T_4535 ? T_3370_bits_data : iofSelReg;
  assign T_4557 = T_3457 == 1'h0;
  assign T_4559 = T_4557 | T_3619_0;
  assign T_4561 = T_3493 == 1'h0;
  assign T_4563 = T_4561 | T_3619_4;
  assign T_4565 = T_3529 == 1'h0;
  assign T_4567 = T_4565 | T_3619_8;
  assign T_4569 = T_3556 == 1'h0;
  assign T_4571 = T_4569 | T_3619_11;
  assign T_4573 = T_3592 == 1'h0;
  assign T_4575 = T_4573 | T_3619_15;
  assign T_4577 = T_3466 == 1'h0;
  assign T_4579 = T_4577 | T_3619_1;
  assign T_4581 = T_3502 == 1'h0;
  assign T_4583 = T_4581 | T_3619_5;
  assign T_4585 = T_3547 == 1'h0;
  assign T_4587 = T_4585 | T_3619_10;
  assign T_4589 = T_3583 == 1'h0;
  assign T_4591 = T_4589 | T_3619_14;
  assign T_4593 = T_3511 == 1'h0;
  assign T_4595 = T_4593 | T_3619_6;
  assign T_4597 = T_3475 == 1'h0;
  assign T_4599 = T_4597 | T_3619_2;
  assign T_4601 = T_3574 == 1'h0;
  assign T_4603 = T_4601 | T_3619_13;
  assign T_4605 = T_3538 == 1'h0;
  assign T_4607 = T_4605 | T_3619_9;
  assign T_4609 = T_3520 == 1'h0;
  assign T_4611 = T_4609 | T_3619_7;
  assign T_4613 = T_3484 == 1'h0;
  assign T_4615 = T_4613 | T_3619_3;
  assign T_4617 = T_3601 == 1'h0;
  assign T_4619 = T_4617 | T_3619_16;
  assign T_4621 = T_3565 == 1'h0;
  assign T_4623 = T_4621 | T_3619_12;
  assign T_4704_0 = T_4559;
  assign T_4704_1 = T_4563;
  assign T_4704_2 = T_4567;
  assign T_4704_3 = T_4571;
  assign T_4704_4 = T_4575;
  assign T_4704_5 = T_4579;
  assign T_4704_6 = T_4583;
  assign T_4704_7 = T_4587;
  assign T_4704_8 = T_4591;
  assign T_4704_9 = T_4595;
  assign T_4704_10 = T_4599;
  assign T_4704_11 = T_4603;
  assign T_4704_12 = T_4607;
  assign T_4704_13 = T_4611;
  assign T_4704_14 = T_4615;
  assign T_4704_15 = T_4619;
  assign T_4704_16 = T_4623;
  assign T_4704_17 = 1'h1;
  assign T_4704_18 = 1'h1;
  assign T_4704_19 = 1'h1;
  assign T_4704_20 = 1'h1;
  assign T_4704_21 = 1'h1;
  assign T_4704_22 = 1'h1;
  assign T_4704_23 = 1'h1;
  assign T_4704_24 = 1'h1;
  assign T_4704_25 = 1'h1;
  assign T_4704_26 = 1'h1;
  assign T_4704_27 = 1'h1;
  assign T_4704_28 = 1'h1;
  assign T_4704_29 = 1'h1;
  assign T_4704_30 = 1'h1;
  assign T_4704_31 = 1'h1;
  assign T_4742 = T_4557 | T_3624_0;
  assign T_4746 = T_4561 | T_3624_4;
  assign T_4750 = T_4565 | T_3624_8;
  assign T_4754 = T_4569 | T_3624_11;
  assign T_4758 = T_4573 | T_3624_15;
  assign T_4762 = T_4577 | T_3624_1;
  assign T_4766 = T_4581 | T_3624_5;
  assign T_4770 = T_4585 | T_3624_10;
  assign T_4774 = T_4589 | T_3624_14;
  assign T_4778 = T_4593 | T_3624_6;
  assign T_4782 = T_4597 | T_3624_2;
  assign T_4786 = T_4601 | T_3624_13;
  assign T_4790 = T_4605 | T_3624_9;
  assign T_4794 = T_4609 | T_3624_7;
  assign T_4798 = T_4613 | T_3624_3;
  assign T_4802 = T_4617 | T_3624_16;
  assign T_4806 = T_4621 | T_3624_12;
  assign T_4887_0 = T_4742;
  assign T_4887_1 = T_4746;
  assign T_4887_2 = T_4750;
  assign T_4887_3 = T_4754;
  assign T_4887_4 = T_4758;
  assign T_4887_5 = T_4762;
  assign T_4887_6 = T_4766;
  assign T_4887_7 = T_4770;
  assign T_4887_8 = T_4774;
  assign T_4887_9 = T_4778;
  assign T_4887_10 = T_4782;
  assign T_4887_11 = T_4786;
  assign T_4887_12 = T_4790;
  assign T_4887_13 = T_4794;
  assign T_4887_14 = T_4798;
  assign T_4887_15 = T_4802;
  assign T_4887_16 = T_4806;
  assign T_4887_17 = 1'h1;
  assign T_4887_18 = 1'h1;
  assign T_4887_19 = 1'h1;
  assign T_4887_20 = 1'h1;
  assign T_4887_21 = 1'h1;
  assign T_4887_22 = 1'h1;
  assign T_4887_23 = 1'h1;
  assign T_4887_24 = 1'h1;
  assign T_4887_25 = 1'h1;
  assign T_4887_26 = 1'h1;
  assign T_4887_27 = 1'h1;
  assign T_4887_28 = 1'h1;
  assign T_4887_29 = 1'h1;
  assign T_4887_30 = 1'h1;
  assign T_4887_31 = 1'h1;
  assign T_4925 = T_4557 | T_3629_0;
  assign T_4929 = T_4561 | T_3629_4;
  assign T_4933 = T_4565 | T_3629_8;
  assign T_4937 = T_4569 | T_3629_11;
  assign T_4941 = T_4573 | T_3629_15;
  assign T_4945 = T_4577 | T_3629_1;
  assign T_4949 = T_4581 | T_3629_5;
  assign T_4953 = T_4585 | T_3629_10;
  assign T_4957 = T_4589 | T_3629_14;
  assign T_4961 = T_4593 | T_3629_6;
  assign T_4965 = T_4597 | T_3629_2;
  assign T_4969 = T_4601 | T_3629_13;
  assign T_4973 = T_4605 | T_3629_9;
  assign T_4977 = T_4609 | T_3629_7;
  assign T_4981 = T_4613 | T_3629_3;
  assign T_4985 = T_4617 | T_3629_16;
  assign T_4989 = T_4621 | T_3629_12;
  assign T_5070_0 = T_4925;
  assign T_5070_1 = T_4929;
  assign T_5070_2 = T_4933;
  assign T_5070_3 = T_4937;
  assign T_5070_4 = T_4941;
  assign T_5070_5 = T_4945;
  assign T_5070_6 = T_4949;
  assign T_5070_7 = T_4953;
  assign T_5070_8 = T_4957;
  assign T_5070_9 = T_4961;
  assign T_5070_10 = T_4965;
  assign T_5070_11 = T_4969;
  assign T_5070_12 = T_4973;
  assign T_5070_13 = T_4977;
  assign T_5070_14 = T_4981;
  assign T_5070_15 = T_4985;
  assign T_5070_16 = T_4989;
  assign T_5070_17 = 1'h1;
  assign T_5070_18 = 1'h1;
  assign T_5070_19 = 1'h1;
  assign T_5070_20 = 1'h1;
  assign T_5070_21 = 1'h1;
  assign T_5070_22 = 1'h1;
  assign T_5070_23 = 1'h1;
  assign T_5070_24 = 1'h1;
  assign T_5070_25 = 1'h1;
  assign T_5070_26 = 1'h1;
  assign T_5070_27 = 1'h1;
  assign T_5070_28 = 1'h1;
  assign T_5070_29 = 1'h1;
  assign T_5070_30 = 1'h1;
  assign T_5070_31 = 1'h1;
  assign T_5108 = T_4557 | T_3634_0;
  assign T_5112 = T_4561 | T_3634_4;
  assign T_5116 = T_4565 | T_3634_8;
  assign T_5120 = T_4569 | T_3634_11;
  assign T_5124 = T_4573 | T_3634_15;
  assign T_5128 = T_4577 | T_3634_1;
  assign T_5132 = T_4581 | T_3634_5;
  assign T_5136 = T_4585 | T_3634_10;
  assign T_5140 = T_4589 | T_3634_14;
  assign T_5144 = T_4593 | T_3634_6;
  assign T_5148 = T_4597 | T_3634_2;
  assign T_5152 = T_4601 | T_3634_13;
  assign T_5156 = T_4605 | T_3634_9;
  assign T_5160 = T_4609 | T_3634_7;
  assign T_5164 = T_4613 | T_3634_3;
  assign T_5168 = T_4617 | T_3634_16;
  assign T_5172 = T_4621 | T_3634_12;
  assign T_5253_0 = T_5108;
  assign T_5253_1 = T_5112;
  assign T_5253_2 = T_5116;
  assign T_5253_3 = T_5120;
  assign T_5253_4 = T_5124;
  assign T_5253_5 = T_5128;
  assign T_5253_6 = T_5132;
  assign T_5253_7 = T_5136;
  assign T_5253_8 = T_5140;
  assign T_5253_9 = T_5144;
  assign T_5253_10 = T_5148;
  assign T_5253_11 = T_5152;
  assign T_5253_12 = T_5156;
  assign T_5253_13 = T_5160;
  assign T_5253_14 = T_5164;
  assign T_5253_15 = T_5168;
  assign T_5253_16 = T_5172;
  assign T_5253_17 = 1'h1;
  assign T_5253_18 = 1'h1;
  assign T_5253_19 = 1'h1;
  assign T_5253_20 = 1'h1;
  assign T_5253_21 = 1'h1;
  assign T_5253_22 = 1'h1;
  assign T_5253_23 = 1'h1;
  assign T_5253_24 = 1'h1;
  assign T_5253_25 = 1'h1;
  assign T_5253_26 = 1'h1;
  assign T_5253_27 = 1'h1;
  assign T_5253_28 = 1'h1;
  assign T_5253_29 = 1'h1;
  assign T_5253_30 = 1'h1;
  assign T_5253_31 = 1'h1;
  assign T_5288 = T_3370_bits_index[0];
  assign T_5289 = T_3370_bits_index[1];
  assign T_5290 = T_3370_bits_index[2];
  assign T_5291 = T_3370_bits_index[3];
  assign T_5292 = T_3370_bits_index[4];
  assign T_5298 = {T_5289,T_5288};
  assign T_5299 = {T_5292,T_5291};
  assign T_5300 = {T_5299,T_5290};
  assign T_5301 = {T_5300,T_5298};
  assign GEN_0 = GEN_45;
  assign GEN_15 = 5'h1 == T_5301 ? T_4704_1 : T_4704_0;
  assign GEN_16 = 5'h2 == T_5301 ? T_4704_2 : GEN_15;
  assign GEN_17 = 5'h3 == T_5301 ? T_4704_3 : GEN_16;
  assign GEN_18 = 5'h4 == T_5301 ? T_4704_4 : GEN_17;
  assign GEN_19 = 5'h5 == T_5301 ? T_4704_5 : GEN_18;
  assign GEN_20 = 5'h6 == T_5301 ? T_4704_6 : GEN_19;
  assign GEN_21 = 5'h7 == T_5301 ? T_4704_7 : GEN_20;
  assign GEN_22 = 5'h8 == T_5301 ? T_4704_8 : GEN_21;
  assign GEN_23 = 5'h9 == T_5301 ? T_4704_9 : GEN_22;
  assign GEN_24 = 5'ha == T_5301 ? T_4704_10 : GEN_23;
  assign GEN_25 = 5'hb == T_5301 ? T_4704_11 : GEN_24;
  assign GEN_26 = 5'hc == T_5301 ? T_4704_12 : GEN_25;
  assign GEN_27 = 5'hd == T_5301 ? T_4704_13 : GEN_26;
  assign GEN_28 = 5'he == T_5301 ? T_4704_14 : GEN_27;
  assign GEN_29 = 5'hf == T_5301 ? T_4704_15 : GEN_28;
  assign GEN_30 = 5'h10 == T_5301 ? T_4704_16 : GEN_29;
  assign GEN_31 = 5'h11 == T_5301 ? T_4704_17 : GEN_30;
  assign GEN_32 = 5'h12 == T_5301 ? T_4704_18 : GEN_31;
  assign GEN_33 = 5'h13 == T_5301 ? T_4704_19 : GEN_32;
  assign GEN_34 = 5'h14 == T_5301 ? T_4704_20 : GEN_33;
  assign GEN_35 = 5'h15 == T_5301 ? T_4704_21 : GEN_34;
  assign GEN_36 = 5'h16 == T_5301 ? T_4704_22 : GEN_35;
  assign GEN_37 = 5'h17 == T_5301 ? T_4704_23 : GEN_36;
  assign GEN_38 = 5'h18 == T_5301 ? T_4704_24 : GEN_37;
  assign GEN_39 = 5'h19 == T_5301 ? T_4704_25 : GEN_38;
  assign GEN_40 = 5'h1a == T_5301 ? T_4704_26 : GEN_39;
  assign GEN_41 = 5'h1b == T_5301 ? T_4704_27 : GEN_40;
  assign GEN_42 = 5'h1c == T_5301 ? T_4704_28 : GEN_41;
  assign GEN_43 = 5'h1d == T_5301 ? T_4704_29 : GEN_42;
  assign GEN_44 = 5'h1e == T_5301 ? T_4704_30 : GEN_43;
  assign GEN_45 = 5'h1f == T_5301 ? T_4704_31 : GEN_44;
  assign GEN_1 = GEN_76;
  assign GEN_46 = 5'h1 == T_5301 ? T_4887_1 : T_4887_0;
  assign GEN_47 = 5'h2 == T_5301 ? T_4887_2 : GEN_46;
  assign GEN_48 = 5'h3 == T_5301 ? T_4887_3 : GEN_47;
  assign GEN_49 = 5'h4 == T_5301 ? T_4887_4 : GEN_48;
  assign GEN_50 = 5'h5 == T_5301 ? T_4887_5 : GEN_49;
  assign GEN_51 = 5'h6 == T_5301 ? T_4887_6 : GEN_50;
  assign GEN_52 = 5'h7 == T_5301 ? T_4887_7 : GEN_51;
  assign GEN_53 = 5'h8 == T_5301 ? T_4887_8 : GEN_52;
  assign GEN_54 = 5'h9 == T_5301 ? T_4887_9 : GEN_53;
  assign GEN_55 = 5'ha == T_5301 ? T_4887_10 : GEN_54;
  assign GEN_56 = 5'hb == T_5301 ? T_4887_11 : GEN_55;
  assign GEN_57 = 5'hc == T_5301 ? T_4887_12 : GEN_56;
  assign GEN_58 = 5'hd == T_5301 ? T_4887_13 : GEN_57;
  assign GEN_59 = 5'he == T_5301 ? T_4887_14 : GEN_58;
  assign GEN_60 = 5'hf == T_5301 ? T_4887_15 : GEN_59;
  assign GEN_61 = 5'h10 == T_5301 ? T_4887_16 : GEN_60;
  assign GEN_62 = 5'h11 == T_5301 ? T_4887_17 : GEN_61;
  assign GEN_63 = 5'h12 == T_5301 ? T_4887_18 : GEN_62;
  assign GEN_64 = 5'h13 == T_5301 ? T_4887_19 : GEN_63;
  assign GEN_65 = 5'h14 == T_5301 ? T_4887_20 : GEN_64;
  assign GEN_66 = 5'h15 == T_5301 ? T_4887_21 : GEN_65;
  assign GEN_67 = 5'h16 == T_5301 ? T_4887_22 : GEN_66;
  assign GEN_68 = 5'h17 == T_5301 ? T_4887_23 : GEN_67;
  assign GEN_69 = 5'h18 == T_5301 ? T_4887_24 : GEN_68;
  assign GEN_70 = 5'h19 == T_5301 ? T_4887_25 : GEN_69;
  assign GEN_71 = 5'h1a == T_5301 ? T_4887_26 : GEN_70;
  assign GEN_72 = 5'h1b == T_5301 ? T_4887_27 : GEN_71;
  assign GEN_73 = 5'h1c == T_5301 ? T_4887_28 : GEN_72;
  assign GEN_74 = 5'h1d == T_5301 ? T_4887_29 : GEN_73;
  assign GEN_75 = 5'h1e == T_5301 ? T_4887_30 : GEN_74;
  assign GEN_76 = 5'h1f == T_5301 ? T_4887_31 : GEN_75;
  assign T_5318 = T_3370_bits_read ? GEN_0 : GEN_1;
  assign GEN_2 = GEN_107;
  assign GEN_77 = 5'h1 == T_5301 ? T_5070_1 : T_5070_0;
  assign GEN_78 = 5'h2 == T_5301 ? T_5070_2 : GEN_77;
  assign GEN_79 = 5'h3 == T_5301 ? T_5070_3 : GEN_78;
  assign GEN_80 = 5'h4 == T_5301 ? T_5070_4 : GEN_79;
  assign GEN_81 = 5'h5 == T_5301 ? T_5070_5 : GEN_80;
  assign GEN_82 = 5'h6 == T_5301 ? T_5070_6 : GEN_81;
  assign GEN_83 = 5'h7 == T_5301 ? T_5070_7 : GEN_82;
  assign GEN_84 = 5'h8 == T_5301 ? T_5070_8 : GEN_83;
  assign GEN_85 = 5'h9 == T_5301 ? T_5070_9 : GEN_84;
  assign GEN_86 = 5'ha == T_5301 ? T_5070_10 : GEN_85;
  assign GEN_87 = 5'hb == T_5301 ? T_5070_11 : GEN_86;
  assign GEN_88 = 5'hc == T_5301 ? T_5070_12 : GEN_87;
  assign GEN_89 = 5'hd == T_5301 ? T_5070_13 : GEN_88;
  assign GEN_90 = 5'he == T_5301 ? T_5070_14 : GEN_89;
  assign GEN_91 = 5'hf == T_5301 ? T_5070_15 : GEN_90;
  assign GEN_92 = 5'h10 == T_5301 ? T_5070_16 : GEN_91;
  assign GEN_93 = 5'h11 == T_5301 ? T_5070_17 : GEN_92;
  assign GEN_94 = 5'h12 == T_5301 ? T_5070_18 : GEN_93;
  assign GEN_95 = 5'h13 == T_5301 ? T_5070_19 : GEN_94;
  assign GEN_96 = 5'h14 == T_5301 ? T_5070_20 : GEN_95;
  assign GEN_97 = 5'h15 == T_5301 ? T_5070_21 : GEN_96;
  assign GEN_98 = 5'h16 == T_5301 ? T_5070_22 : GEN_97;
  assign GEN_99 = 5'h17 == T_5301 ? T_5070_23 : GEN_98;
  assign GEN_100 = 5'h18 == T_5301 ? T_5070_24 : GEN_99;
  assign GEN_101 = 5'h19 == T_5301 ? T_5070_25 : GEN_100;
  assign GEN_102 = 5'h1a == T_5301 ? T_5070_26 : GEN_101;
  assign GEN_103 = 5'h1b == T_5301 ? T_5070_27 : GEN_102;
  assign GEN_104 = 5'h1c == T_5301 ? T_5070_28 : GEN_103;
  assign GEN_105 = 5'h1d == T_5301 ? T_5070_29 : GEN_104;
  assign GEN_106 = 5'h1e == T_5301 ? T_5070_30 : GEN_105;
  assign GEN_107 = 5'h1f == T_5301 ? T_5070_31 : GEN_106;
  assign GEN_3 = GEN_138;
  assign GEN_108 = 5'h1 == T_5301 ? T_5253_1 : T_5253_0;
  assign GEN_109 = 5'h2 == T_5301 ? T_5253_2 : GEN_108;
  assign GEN_110 = 5'h3 == T_5301 ? T_5253_3 : GEN_109;
  assign GEN_111 = 5'h4 == T_5301 ? T_5253_4 : GEN_110;
  assign GEN_112 = 5'h5 == T_5301 ? T_5253_5 : GEN_111;
  assign GEN_113 = 5'h6 == T_5301 ? T_5253_6 : GEN_112;
  assign GEN_114 = 5'h7 == T_5301 ? T_5253_7 : GEN_113;
  assign GEN_115 = 5'h8 == T_5301 ? T_5253_8 : GEN_114;
  assign GEN_116 = 5'h9 == T_5301 ? T_5253_9 : GEN_115;
  assign GEN_117 = 5'ha == T_5301 ? T_5253_10 : GEN_116;
  assign GEN_118 = 5'hb == T_5301 ? T_5253_11 : GEN_117;
  assign GEN_119 = 5'hc == T_5301 ? T_5253_12 : GEN_118;
  assign GEN_120 = 5'hd == T_5301 ? T_5253_13 : GEN_119;
  assign GEN_121 = 5'he == T_5301 ? T_5253_14 : GEN_120;
  assign GEN_122 = 5'hf == T_5301 ? T_5253_15 : GEN_121;
  assign GEN_123 = 5'h10 == T_5301 ? T_5253_16 : GEN_122;
  assign GEN_124 = 5'h11 == T_5301 ? T_5253_17 : GEN_123;
  assign GEN_125 = 5'h12 == T_5301 ? T_5253_18 : GEN_124;
  assign GEN_126 = 5'h13 == T_5301 ? T_5253_19 : GEN_125;
  assign GEN_127 = 5'h14 == T_5301 ? T_5253_20 : GEN_126;
  assign GEN_128 = 5'h15 == T_5301 ? T_5253_21 : GEN_127;
  assign GEN_129 = 5'h16 == T_5301 ? T_5253_22 : GEN_128;
  assign GEN_130 = 5'h17 == T_5301 ? T_5253_23 : GEN_129;
  assign GEN_131 = 5'h18 == T_5301 ? T_5253_24 : GEN_130;
  assign GEN_132 = 5'h19 == T_5301 ? T_5253_25 : GEN_131;
  assign GEN_133 = 5'h1a == T_5301 ? T_5253_26 : GEN_132;
  assign GEN_134 = 5'h1b == T_5301 ? T_5253_27 : GEN_133;
  assign GEN_135 = 5'h1c == T_5301 ? T_5253_28 : GEN_134;
  assign GEN_136 = 5'h1d == T_5301 ? T_5253_29 : GEN_135;
  assign GEN_137 = 5'h1e == T_5301 ? T_5253_30 : GEN_136;
  assign GEN_138 = 5'h1f == T_5301 ? T_5253_31 : GEN_137;
  assign T_5321 = T_3370_bits_read ? GEN_2 : GEN_3;
  assign T_5322 = T_3370_ready & T_5318;
  assign T_5323 = T_3295_valid & T_5318;
  assign T_5324 = T_3334_ready & T_5321;
  assign T_5325 = T_3370_valid & T_5321;
  assign T_5327 = 32'h1 << T_5301;
  assign T_5328 = {T_3493,T_3457};
  assign T_5329 = {T_3556,T_3529};
  assign T_5330 = {T_5329,T_5328};
  assign T_5331 = {T_3466,T_3592};
  assign T_5332 = {T_3547,T_3502};
  assign T_5333 = {T_5332,T_5331};
  assign T_5334 = {T_5333,T_5330};
  assign T_5335 = {T_3511,T_3583};
  assign T_5336 = {T_3574,T_3475};
  assign T_5337 = {T_5336,T_5335};
  assign T_5338 = {T_3520,T_3538};
  assign T_5339 = {T_3601,T_3484};
  assign T_5340 = {T_5339,T_5338};
  assign T_5341 = {T_5340,T_5337};
  assign T_5342 = {T_5341,T_5334};
  assign T_5343 = {1'h1,T_3565};
  assign T_5345 = {2'h3,T_5343};
  assign T_5349 = {4'hf,T_5345};
  assign T_5357 = {8'hff,T_5349};
  assign T_5358 = {T_5357,T_5342};
  assign T_5359 = T_5327 & T_5358;
  assign T_5394 = T_3295_valid & T_3370_ready;
  assign T_5395 = T_5394 & T_3370_bits_read;
  assign T_5396 = T_5359[0];
  assign T_5397 = T_5395 & T_5396;
  assign T_5400 = T_3370_bits_read == 1'h0;
  assign T_5401 = T_5394 & T_5400;
  assign T_5403 = T_5401 & T_5396;
  assign T_5404 = T_3370_valid & T_3334_ready;
  assign T_5405 = T_5404 & T_3370_bits_read;
  assign T_5407 = T_5405 & T_5396;
  assign T_5411 = T_5404 & T_5400;
  assign T_5413 = T_5411 & T_5396;
  assign T_5416 = T_5359[1];
  assign T_5417 = T_5395 & T_5416;
  assign T_5423 = T_5401 & T_5416;
  assign T_5427 = T_5405 & T_5416;
  assign T_5433 = T_5411 & T_5416;
  assign T_5436 = T_5359[2];
  assign T_5437 = T_5395 & T_5436;
  assign T_5443 = T_5401 & T_5436;
  assign T_5447 = T_5405 & T_5436;
  assign T_5453 = T_5411 & T_5436;
  assign T_5456 = T_5359[3];
  assign T_5457 = T_5395 & T_5456;
  assign T_5463 = T_5401 & T_5456;
  assign T_5467 = T_5405 & T_5456;
  assign T_5473 = T_5411 & T_5456;
  assign T_5476 = T_5359[4];
  assign T_5477 = T_5395 & T_5476;
  assign T_5483 = T_5401 & T_5476;
  assign T_5487 = T_5405 & T_5476;
  assign T_5493 = T_5411 & T_5476;
  assign T_5496 = T_5359[5];
  assign T_5497 = T_5395 & T_5496;
  assign T_5503 = T_5401 & T_5496;
  assign T_5507 = T_5405 & T_5496;
  assign T_5513 = T_5411 & T_5496;
  assign T_5516 = T_5359[6];
  assign T_5517 = T_5395 & T_5516;
  assign T_5523 = T_5401 & T_5516;
  assign T_5527 = T_5405 & T_5516;
  assign T_5533 = T_5411 & T_5516;
  assign T_5536 = T_5359[7];
  assign T_5537 = T_5395 & T_5536;
  assign T_5543 = T_5401 & T_5536;
  assign T_5547 = T_5405 & T_5536;
  assign T_5553 = T_5411 & T_5536;
  assign T_5556 = T_5359[8];
  assign T_5557 = T_5395 & T_5556;
  assign T_5563 = T_5401 & T_5556;
  assign T_5567 = T_5405 & T_5556;
  assign T_5573 = T_5411 & T_5556;
  assign T_5576 = T_5359[9];
  assign T_5577 = T_5395 & T_5576;
  assign T_5583 = T_5401 & T_5576;
  assign T_5587 = T_5405 & T_5576;
  assign T_5593 = T_5411 & T_5576;
  assign T_5596 = T_5359[10];
  assign T_5597 = T_5395 & T_5596;
  assign T_5603 = T_5401 & T_5596;
  assign T_5607 = T_5405 & T_5596;
  assign T_5613 = T_5411 & T_5596;
  assign T_5616 = T_5359[11];
  assign T_5617 = T_5395 & T_5616;
  assign T_5623 = T_5401 & T_5616;
  assign T_5627 = T_5405 & T_5616;
  assign T_5633 = T_5411 & T_5616;
  assign T_5636 = T_5359[12];
  assign T_5637 = T_5395 & T_5636;
  assign T_5643 = T_5401 & T_5636;
  assign T_5647 = T_5405 & T_5636;
  assign T_5653 = T_5411 & T_5636;
  assign T_5656 = T_5359[13];
  assign T_5657 = T_5395 & T_5656;
  assign T_5663 = T_5401 & T_5656;
  assign T_5667 = T_5405 & T_5656;
  assign T_5673 = T_5411 & T_5656;
  assign T_5676 = T_5359[14];
  assign T_5677 = T_5395 & T_5676;
  assign T_5683 = T_5401 & T_5676;
  assign T_5687 = T_5405 & T_5676;
  assign T_5693 = T_5411 & T_5676;
  assign T_5696 = T_5359[15];
  assign T_5697 = T_5395 & T_5696;
  assign T_5703 = T_5401 & T_5696;
  assign T_5707 = T_5405 & T_5696;
  assign T_5713 = T_5411 & T_5696;
  assign T_5716 = T_5359[16];
  assign T_5717 = T_5395 & T_5716;
  assign T_5723 = T_5401 & T_5716;
  assign T_5727 = T_5405 & T_5716;
  assign T_5733 = T_5411 & T_5716;
  assign T_6137_0 = T_3457;
  assign T_6137_1 = T_3493;
  assign T_6137_2 = T_3529;
  assign T_6137_3 = T_3556;
  assign T_6137_4 = T_3592;
  assign T_6137_5 = T_3466;
  assign T_6137_6 = T_3502;
  assign T_6137_7 = T_3547;
  assign T_6137_8 = T_3583;
  assign T_6137_9 = T_3511;
  assign T_6137_10 = T_3475;
  assign T_6137_11 = T_3574;
  assign T_6137_12 = T_3538;
  assign T_6137_13 = T_3520;
  assign T_6137_14 = T_3484;
  assign T_6137_15 = T_3601;
  assign T_6137_16 = T_3565;
  assign T_6137_17 = 1'h1;
  assign T_6137_18 = 1'h1;
  assign T_6137_19 = 1'h1;
  assign T_6137_20 = 1'h1;
  assign T_6137_21 = 1'h1;
  assign T_6137_22 = 1'h1;
  assign T_6137_23 = 1'h1;
  assign T_6137_24 = 1'h1;
  assign T_6137_25 = 1'h1;
  assign T_6137_26 = 1'h1;
  assign T_6137_27 = 1'h1;
  assign T_6137_28 = 1'h1;
  assign T_6137_29 = 1'h1;
  assign T_6137_30 = 1'h1;
  assign T_6137_31 = 1'h1;
  assign T_6208_0 = valueReg;
  assign T_6208_1 = T_4047;
  assign T_6208_2 = T_4219;
  assign T_6208_3 = portReg;
  assign T_6208_4 = T_4511;
  assign T_6208_5 = dsReg;
  assign T_6208_6 = riseIeReg;
  assign T_6208_7 = riseIpReg;
  assign T_6208_8 = fallIeReg;
  assign T_6208_9 = fallIpReg;
  assign T_6208_10 = highIeReg;
  assign T_6208_11 = highIpReg;
  assign T_6208_12 = lowIeReg;
  assign T_6208_13 = lowIpReg;
  assign T_6208_14 = T_4007;
  assign T_6208_15 = iofSelReg;
  assign T_6208_16 = xorReg;
  assign T_6208_17 = 32'h0;
  assign T_6208_18 = 32'h0;
  assign T_6208_19 = 32'h0;
  assign T_6208_20 = 32'h0;
  assign T_6208_21 = 32'h0;
  assign T_6208_22 = 32'h0;
  assign T_6208_23 = 32'h0;
  assign T_6208_24 = 32'h0;
  assign T_6208_25 = 32'h0;
  assign T_6208_26 = 32'h0;
  assign T_6208_27 = 32'h0;
  assign T_6208_28 = 32'h0;
  assign T_6208_29 = 32'h0;
  assign T_6208_30 = 32'h0;
  assign T_6208_31 = 32'h0;
  assign GEN_4 = GEN_169;
  assign GEN_139 = 5'h1 == T_5301 ? T_6137_1 : T_6137_0;
  assign GEN_140 = 5'h2 == T_5301 ? T_6137_2 : GEN_139;
  assign GEN_141 = 5'h3 == T_5301 ? T_6137_3 : GEN_140;
  assign GEN_142 = 5'h4 == T_5301 ? T_6137_4 : GEN_141;
  assign GEN_143 = 5'h5 == T_5301 ? T_6137_5 : GEN_142;
  assign GEN_144 = 5'h6 == T_5301 ? T_6137_6 : GEN_143;
  assign GEN_145 = 5'h7 == T_5301 ? T_6137_7 : GEN_144;
  assign GEN_146 = 5'h8 == T_5301 ? T_6137_8 : GEN_145;
  assign GEN_147 = 5'h9 == T_5301 ? T_6137_9 : GEN_146;
  assign GEN_148 = 5'ha == T_5301 ? T_6137_10 : GEN_147;
  assign GEN_149 = 5'hb == T_5301 ? T_6137_11 : GEN_148;
  assign GEN_150 = 5'hc == T_5301 ? T_6137_12 : GEN_149;
  assign GEN_151 = 5'hd == T_5301 ? T_6137_13 : GEN_150;
  assign GEN_152 = 5'he == T_5301 ? T_6137_14 : GEN_151;
  assign GEN_153 = 5'hf == T_5301 ? T_6137_15 : GEN_152;
  assign GEN_154 = 5'h10 == T_5301 ? T_6137_16 : GEN_153;
  assign GEN_155 = 5'h11 == T_5301 ? T_6137_17 : GEN_154;
  assign GEN_156 = 5'h12 == T_5301 ? T_6137_18 : GEN_155;
  assign GEN_157 = 5'h13 == T_5301 ? T_6137_19 : GEN_156;
  assign GEN_158 = 5'h14 == T_5301 ? T_6137_20 : GEN_157;
  assign GEN_159 = 5'h15 == T_5301 ? T_6137_21 : GEN_158;
  assign GEN_160 = 5'h16 == T_5301 ? T_6137_22 : GEN_159;
  assign GEN_161 = 5'h17 == T_5301 ? T_6137_23 : GEN_160;
  assign GEN_162 = 5'h18 == T_5301 ? T_6137_24 : GEN_161;
  assign GEN_163 = 5'h19 == T_5301 ? T_6137_25 : GEN_162;
  assign GEN_164 = 5'h1a == T_5301 ? T_6137_26 : GEN_163;
  assign GEN_165 = 5'h1b == T_5301 ? T_6137_27 : GEN_164;
  assign GEN_166 = 5'h1c == T_5301 ? T_6137_28 : GEN_165;
  assign GEN_167 = 5'h1d == T_5301 ? T_6137_29 : GEN_166;
  assign GEN_168 = 5'h1e == T_5301 ? T_6137_30 : GEN_167;
  assign GEN_169 = 5'h1f == T_5301 ? T_6137_31 : GEN_168;
  assign GEN_5 = GEN_200;
  assign GEN_170 = 5'h1 == T_5301 ? T_6208_1 : T_6208_0;
  assign GEN_171 = 5'h2 == T_5301 ? T_6208_2 : GEN_170;
  assign GEN_172 = 5'h3 == T_5301 ? T_6208_3 : GEN_171;
  assign GEN_173 = 5'h4 == T_5301 ? T_6208_4 : GEN_172;
  assign GEN_174 = 5'h5 == T_5301 ? T_6208_5 : GEN_173;
  assign GEN_175 = 5'h6 == T_5301 ? T_6208_6 : GEN_174;
  assign GEN_176 = 5'h7 == T_5301 ? T_6208_7 : GEN_175;
  assign GEN_177 = 5'h8 == T_5301 ? T_6208_8 : GEN_176;
  assign GEN_178 = 5'h9 == T_5301 ? T_6208_9 : GEN_177;
  assign GEN_179 = 5'ha == T_5301 ? T_6208_10 : GEN_178;
  assign GEN_180 = 5'hb == T_5301 ? T_6208_11 : GEN_179;
  assign GEN_181 = 5'hc == T_5301 ? T_6208_12 : GEN_180;
  assign GEN_182 = 5'hd == T_5301 ? T_6208_13 : GEN_181;
  assign GEN_183 = 5'he == T_5301 ? T_6208_14 : GEN_182;
  assign GEN_184 = 5'hf == T_5301 ? T_6208_15 : GEN_183;
  assign GEN_185 = 5'h10 == T_5301 ? T_6208_16 : GEN_184;
  assign GEN_186 = 5'h11 == T_5301 ? T_6208_17 : GEN_185;
  assign GEN_187 = 5'h12 == T_5301 ? T_6208_18 : GEN_186;
  assign GEN_188 = 5'h13 == T_5301 ? T_6208_19 : GEN_187;
  assign GEN_189 = 5'h14 == T_5301 ? T_6208_20 : GEN_188;
  assign GEN_190 = 5'h15 == T_5301 ? T_6208_21 : GEN_189;
  assign GEN_191 = 5'h16 == T_5301 ? T_6208_22 : GEN_190;
  assign GEN_192 = 5'h17 == T_5301 ? T_6208_23 : GEN_191;
  assign GEN_193 = 5'h18 == T_5301 ? T_6208_24 : GEN_192;
  assign GEN_194 = 5'h19 == T_5301 ? T_6208_25 : GEN_193;
  assign GEN_195 = 5'h1a == T_5301 ? T_6208_26 : GEN_194;
  assign GEN_196 = 5'h1b == T_5301 ? T_6208_27 : GEN_195;
  assign GEN_197 = 5'h1c == T_5301 ? T_6208_28 : GEN_196;
  assign GEN_198 = 5'h1d == T_5301 ? T_6208_29 : GEN_197;
  assign GEN_199 = 5'h1e == T_5301 ? T_6208_30 : GEN_198;
  assign GEN_200 = 5'h1f == T_5301 ? T_6208_31 : GEN_199;
  assign T_6245 = GEN_4 ? GEN_5 : 32'h0;
  assign T_6246 = T_3334_bits_extra[9:8];
  assign T_6248 = T_3334_bits_extra[7:3];
  assign T_6249 = T_3334_bits_extra[2:0];
  assign T_6260_opcode = 3'h0;
  assign T_6260_param = 2'h0;
  assign T_6260_size = T_6249;
  assign T_6260_source = T_6248;
  assign T_6260_sink = 1'h0;
  assign T_6260_addr_lo = T_6246;
  assign T_6260_data = 32'h0;
  assign T_6260_error = 1'h0;
  assign swPinCtrl_0_oval = T_7570;
  assign swPinCtrl_0_oe = T_7571;
  assign swPinCtrl_0_ie = T_7573;
  assign swPinCtrl_0_pue = T_7569;
  assign swPinCtrl_0_ds = T_7572;
  assign swPinCtrl_1_oval = T_7606;
  assign swPinCtrl_1_oe = T_7607;
  assign swPinCtrl_1_ie = T_7609;
  assign swPinCtrl_1_pue = T_7605;
  assign swPinCtrl_1_ds = T_7608;
  assign swPinCtrl_2_oval = T_7642;
  assign swPinCtrl_2_oe = T_7643;
  assign swPinCtrl_2_ie = T_7645;
  assign swPinCtrl_2_pue = T_7641;
  assign swPinCtrl_2_ds = T_7644;
  assign swPinCtrl_3_oval = T_7678;
  assign swPinCtrl_3_oe = T_7679;
  assign swPinCtrl_3_ie = T_7681;
  assign swPinCtrl_3_pue = T_7677;
  assign swPinCtrl_3_ds = T_7680;
  assign swPinCtrl_4_oval = T_7714;
  assign swPinCtrl_4_oe = T_7715;
  assign swPinCtrl_4_ie = T_7717;
  assign swPinCtrl_4_pue = T_7713;
  assign swPinCtrl_4_ds = T_7716;
  assign swPinCtrl_5_oval = T_7750;
  assign swPinCtrl_5_oe = T_7751;
  assign swPinCtrl_5_ie = T_7753;
  assign swPinCtrl_5_pue = T_7749;
  assign swPinCtrl_5_ds = T_7752;
  assign swPinCtrl_6_oval = T_7786;
  assign swPinCtrl_6_oe = T_7787;
  assign swPinCtrl_6_ie = T_7789;
  assign swPinCtrl_6_pue = T_7785;
  assign swPinCtrl_6_ds = T_7788;
  assign swPinCtrl_7_oval = T_7822;
  assign swPinCtrl_7_oe = T_7823;
  assign swPinCtrl_7_ie = T_7825;
  assign swPinCtrl_7_pue = T_7821;
  assign swPinCtrl_7_ds = T_7824;
  assign swPinCtrl_8_oval = T_7858;
  assign swPinCtrl_8_oe = T_7859;
  assign swPinCtrl_8_ie = T_7861;
  assign swPinCtrl_8_pue = T_7857;
  assign swPinCtrl_8_ds = T_7860;
  assign swPinCtrl_9_oval = T_7894;
  assign swPinCtrl_9_oe = T_7895;
  assign swPinCtrl_9_ie = T_7897;
  assign swPinCtrl_9_pue = T_7893;
  assign swPinCtrl_9_ds = T_7896;
  assign swPinCtrl_10_oval = T_7930;
  assign swPinCtrl_10_oe = T_7931;
  assign swPinCtrl_10_ie = T_7933;
  assign swPinCtrl_10_pue = T_7929;
  assign swPinCtrl_10_ds = T_7932;
  assign swPinCtrl_11_oval = T_7966;
  assign swPinCtrl_11_oe = T_7967;
  assign swPinCtrl_11_ie = T_7969;
  assign swPinCtrl_11_pue = T_7965;
  assign swPinCtrl_11_ds = T_7968;
  assign swPinCtrl_12_oval = T_8002;
  assign swPinCtrl_12_oe = T_8003;
  assign swPinCtrl_12_ie = T_8005;
  assign swPinCtrl_12_pue = T_8001;
  assign swPinCtrl_12_ds = T_8004;
  assign swPinCtrl_13_oval = T_8038;
  assign swPinCtrl_13_oe = T_8039;
  assign swPinCtrl_13_ie = T_8041;
  assign swPinCtrl_13_pue = T_8037;
  assign swPinCtrl_13_ds = T_8040;
  assign swPinCtrl_14_oval = T_8074;
  assign swPinCtrl_14_oe = T_8075;
  assign swPinCtrl_14_ie = T_8077;
  assign swPinCtrl_14_pue = T_8073;
  assign swPinCtrl_14_ds = T_8076;
  assign swPinCtrl_15_oval = T_8110;
  assign swPinCtrl_15_oe = T_8111;
  assign swPinCtrl_15_ie = T_8113;
  assign swPinCtrl_15_pue = T_8109;
  assign swPinCtrl_15_ds = T_8112;
  assign swPinCtrl_16_oval = T_8146;
  assign swPinCtrl_16_oe = T_8147;
  assign swPinCtrl_16_ie = T_8149;
  assign swPinCtrl_16_pue = T_8145;
  assign swPinCtrl_16_ds = T_8148;
  assign swPinCtrl_17_oval = T_8182;
  assign swPinCtrl_17_oe = T_8183;
  assign swPinCtrl_17_ie = T_8185;
  assign swPinCtrl_17_pue = T_8181;
  assign swPinCtrl_17_ds = T_8184;
  assign swPinCtrl_18_oval = T_8218;
  assign swPinCtrl_18_oe = T_8219;
  assign swPinCtrl_18_ie = T_8221;
  assign swPinCtrl_18_pue = T_8217;
  assign swPinCtrl_18_ds = T_8220;
  assign swPinCtrl_19_oval = T_8254;
  assign swPinCtrl_19_oe = T_8255;
  assign swPinCtrl_19_ie = T_8257;
  assign swPinCtrl_19_pue = T_8253;
  assign swPinCtrl_19_ds = T_8256;
  assign swPinCtrl_20_oval = T_8290;
  assign swPinCtrl_20_oe = T_8291;
  assign swPinCtrl_20_ie = T_8293;
  assign swPinCtrl_20_pue = T_8289;
  assign swPinCtrl_20_ds = T_8292;
  assign swPinCtrl_21_oval = T_8326;
  assign swPinCtrl_21_oe = T_8327;
  assign swPinCtrl_21_ie = T_8329;
  assign swPinCtrl_21_pue = T_8325;
  assign swPinCtrl_21_ds = T_8328;
  assign swPinCtrl_22_oval = T_8362;
  assign swPinCtrl_22_oe = T_8363;
  assign swPinCtrl_22_ie = T_8365;
  assign swPinCtrl_22_pue = T_8361;
  assign swPinCtrl_22_ds = T_8364;
  assign swPinCtrl_23_oval = T_8398;
  assign swPinCtrl_23_oe = T_8399;
  assign swPinCtrl_23_ie = T_8401;
  assign swPinCtrl_23_pue = T_8397;
  assign swPinCtrl_23_ds = T_8400;
  assign swPinCtrl_24_oval = T_8434;
  assign swPinCtrl_24_oe = T_8435;
  assign swPinCtrl_24_ie = T_8437;
  assign swPinCtrl_24_pue = T_8433;
  assign swPinCtrl_24_ds = T_8436;
  assign swPinCtrl_25_oval = T_8470;
  assign swPinCtrl_25_oe = T_8471;
  assign swPinCtrl_25_ie = T_8473;
  assign swPinCtrl_25_pue = T_8469;
  assign swPinCtrl_25_ds = T_8472;
  assign swPinCtrl_26_oval = T_8506;
  assign swPinCtrl_26_oe = T_8507;
  assign swPinCtrl_26_ie = T_8509;
  assign swPinCtrl_26_pue = T_8505;
  assign swPinCtrl_26_ds = T_8508;
  assign swPinCtrl_27_oval = T_8542;
  assign swPinCtrl_27_oe = T_8543;
  assign swPinCtrl_27_ie = T_8545;
  assign swPinCtrl_27_pue = T_8541;
  assign swPinCtrl_27_ds = T_8544;
  assign swPinCtrl_28_oval = T_8578;
  assign swPinCtrl_28_oe = T_8579;
  assign swPinCtrl_28_ie = T_8581;
  assign swPinCtrl_28_pue = T_8577;
  assign swPinCtrl_28_ds = T_8580;
  assign swPinCtrl_29_oval = T_8614;
  assign swPinCtrl_29_oe = T_8615;
  assign swPinCtrl_29_ie = T_8617;
  assign swPinCtrl_29_pue = T_8613;
  assign swPinCtrl_29_ds = T_8616;
  assign swPinCtrl_30_oval = T_8650;
  assign swPinCtrl_30_oe = T_8651;
  assign swPinCtrl_30_ie = T_8653;
  assign swPinCtrl_30_pue = T_8649;
  assign swPinCtrl_30_ds = T_8652;
  assign swPinCtrl_31_oval = T_8686;
  assign swPinCtrl_31_oe = T_8687;
  assign swPinCtrl_31_ie = T_8689;
  assign swPinCtrl_31_pue = T_8685;
  assign swPinCtrl_31_ds = T_8688;
  assign iof0Ctrl_0_oval = GEN_201;
  assign iof0Ctrl_0_oe = GEN_202;
  assign iof0Ctrl_0_ie = GEN_203;
  assign iof0Ctrl_1_oval = GEN_207;
  assign iof0Ctrl_1_oe = GEN_208;
  assign iof0Ctrl_1_ie = GEN_209;
  assign iof0Ctrl_2_oval = GEN_213;
  assign iof0Ctrl_2_oe = GEN_214;
  assign iof0Ctrl_2_ie = GEN_215;
  assign iof0Ctrl_3_oval = GEN_219;
  assign iof0Ctrl_3_oe = GEN_220;
  assign iof0Ctrl_3_ie = GEN_221;
  assign iof0Ctrl_4_oval = GEN_225;
  assign iof0Ctrl_4_oe = GEN_226;
  assign iof0Ctrl_4_ie = GEN_227;
  assign iof0Ctrl_5_oval = GEN_231;
  assign iof0Ctrl_5_oe = GEN_232;
  assign iof0Ctrl_5_ie = GEN_233;
  assign iof0Ctrl_6_oval = GEN_237;
  assign iof0Ctrl_6_oe = GEN_238;
  assign iof0Ctrl_6_ie = GEN_239;
  assign iof0Ctrl_7_oval = GEN_243;
  assign iof0Ctrl_7_oe = GEN_244;
  assign iof0Ctrl_7_ie = GEN_245;
  assign iof0Ctrl_8_oval = GEN_249;
  assign iof0Ctrl_8_oe = GEN_250;
  assign iof0Ctrl_8_ie = GEN_251;
  assign iof0Ctrl_9_oval = GEN_255;
  assign iof0Ctrl_9_oe = GEN_256;
  assign iof0Ctrl_9_ie = GEN_257;
  assign iof0Ctrl_10_oval = GEN_261;
  assign iof0Ctrl_10_oe = GEN_262;
  assign iof0Ctrl_10_ie = GEN_263;
  assign iof0Ctrl_11_oval = GEN_267;
  assign iof0Ctrl_11_oe = GEN_268;
  assign iof0Ctrl_11_ie = GEN_269;
  assign iof0Ctrl_12_oval = GEN_273;
  assign iof0Ctrl_12_oe = GEN_274;
  assign iof0Ctrl_12_ie = GEN_275;
  assign iof0Ctrl_13_oval = GEN_279;
  assign iof0Ctrl_13_oe = GEN_280;
  assign iof0Ctrl_13_ie = GEN_281;
  assign iof0Ctrl_14_oval = GEN_285;
  assign iof0Ctrl_14_oe = GEN_286;
  assign iof0Ctrl_14_ie = GEN_287;
  assign iof0Ctrl_15_oval = GEN_291;
  assign iof0Ctrl_15_oe = GEN_292;
  assign iof0Ctrl_15_ie = GEN_293;
  assign iof0Ctrl_16_oval = GEN_297;
  assign iof0Ctrl_16_oe = GEN_298;
  assign iof0Ctrl_16_ie = GEN_299;
  assign iof0Ctrl_17_oval = GEN_303;
  assign iof0Ctrl_17_oe = GEN_304;
  assign iof0Ctrl_17_ie = GEN_305;
  assign iof0Ctrl_18_oval = GEN_309;
  assign iof0Ctrl_18_oe = GEN_310;
  assign iof0Ctrl_18_ie = GEN_311;
  assign iof0Ctrl_19_oval = GEN_315;
  assign iof0Ctrl_19_oe = GEN_316;
  assign iof0Ctrl_19_ie = GEN_317;
  assign iof0Ctrl_20_oval = GEN_321;
  assign iof0Ctrl_20_oe = GEN_322;
  assign iof0Ctrl_20_ie = GEN_323;
  assign iof0Ctrl_21_oval = GEN_327;
  assign iof0Ctrl_21_oe = GEN_328;
  assign iof0Ctrl_21_ie = GEN_329;
  assign iof0Ctrl_22_oval = GEN_333;
  assign iof0Ctrl_22_oe = GEN_334;
  assign iof0Ctrl_22_ie = GEN_335;
  assign iof0Ctrl_23_oval = GEN_339;
  assign iof0Ctrl_23_oe = GEN_340;
  assign iof0Ctrl_23_ie = GEN_341;
  assign iof0Ctrl_24_oval = GEN_345;
  assign iof0Ctrl_24_oe = GEN_346;
  assign iof0Ctrl_24_ie = GEN_347;
  assign iof0Ctrl_25_oval = GEN_351;
  assign iof0Ctrl_25_oe = GEN_352;
  assign iof0Ctrl_25_ie = GEN_353;
  assign iof0Ctrl_26_oval = GEN_357;
  assign iof0Ctrl_26_oe = GEN_358;
  assign iof0Ctrl_26_ie = GEN_359;
  assign iof0Ctrl_27_oval = GEN_363;
  assign iof0Ctrl_27_oe = GEN_364;
  assign iof0Ctrl_27_ie = GEN_365;
  assign iof0Ctrl_28_oval = GEN_369;
  assign iof0Ctrl_28_oe = GEN_370;
  assign iof0Ctrl_28_ie = GEN_371;
  assign iof0Ctrl_29_oval = GEN_375;
  assign iof0Ctrl_29_oe = GEN_376;
  assign iof0Ctrl_29_ie = GEN_377;
  assign iof0Ctrl_30_oval = GEN_381;
  assign iof0Ctrl_30_oe = GEN_382;
  assign iof0Ctrl_30_ie = GEN_383;
  assign iof0Ctrl_31_oval = GEN_387;
  assign iof0Ctrl_31_oe = GEN_388;
  assign iof0Ctrl_31_ie = GEN_389;
  assign iof1Ctrl_0_oval = GEN_204;
  assign iof1Ctrl_0_oe = GEN_205;
  assign iof1Ctrl_0_ie = GEN_206;
  assign iof1Ctrl_1_oval = GEN_210;
  assign iof1Ctrl_1_oe = GEN_211;
  assign iof1Ctrl_1_ie = GEN_212;
  assign iof1Ctrl_2_oval = GEN_216;
  assign iof1Ctrl_2_oe = GEN_217;
  assign iof1Ctrl_2_ie = GEN_218;
  assign iof1Ctrl_3_oval = GEN_222;
  assign iof1Ctrl_3_oe = GEN_223;
  assign iof1Ctrl_3_ie = GEN_224;
  assign iof1Ctrl_4_oval = GEN_228;
  assign iof1Ctrl_4_oe = GEN_229;
  assign iof1Ctrl_4_ie = GEN_230;
  assign iof1Ctrl_5_oval = GEN_234;
  assign iof1Ctrl_5_oe = GEN_235;
  assign iof1Ctrl_5_ie = GEN_236;
  assign iof1Ctrl_6_oval = GEN_240;
  assign iof1Ctrl_6_oe = GEN_241;
  assign iof1Ctrl_6_ie = GEN_242;
  assign iof1Ctrl_7_oval = GEN_246;
  assign iof1Ctrl_7_oe = GEN_247;
  assign iof1Ctrl_7_ie = GEN_248;
  assign iof1Ctrl_8_oval = GEN_252;
  assign iof1Ctrl_8_oe = GEN_253;
  assign iof1Ctrl_8_ie = GEN_254;
  assign iof1Ctrl_9_oval = GEN_258;
  assign iof1Ctrl_9_oe = GEN_259;
  assign iof1Ctrl_9_ie = GEN_260;
  assign iof1Ctrl_10_oval = GEN_264;
  assign iof1Ctrl_10_oe = GEN_265;
  assign iof1Ctrl_10_ie = GEN_266;
  assign iof1Ctrl_11_oval = GEN_270;
  assign iof1Ctrl_11_oe = GEN_271;
  assign iof1Ctrl_11_ie = GEN_272;
  assign iof1Ctrl_12_oval = GEN_276;
  assign iof1Ctrl_12_oe = GEN_277;
  assign iof1Ctrl_12_ie = GEN_278;
  assign iof1Ctrl_13_oval = GEN_282;
  assign iof1Ctrl_13_oe = GEN_283;
  assign iof1Ctrl_13_ie = GEN_284;
  assign iof1Ctrl_14_oval = GEN_288;
  assign iof1Ctrl_14_oe = GEN_289;
  assign iof1Ctrl_14_ie = GEN_290;
  assign iof1Ctrl_15_oval = GEN_294;
  assign iof1Ctrl_15_oe = GEN_295;
  assign iof1Ctrl_15_ie = GEN_296;
  assign iof1Ctrl_16_oval = GEN_300;
  assign iof1Ctrl_16_oe = GEN_301;
  assign iof1Ctrl_16_ie = GEN_302;
  assign iof1Ctrl_17_oval = GEN_306;
  assign iof1Ctrl_17_oe = GEN_307;
  assign iof1Ctrl_17_ie = GEN_308;
  assign iof1Ctrl_18_oval = GEN_312;
  assign iof1Ctrl_18_oe = GEN_313;
  assign iof1Ctrl_18_ie = GEN_314;
  assign iof1Ctrl_19_oval = GEN_318;
  assign iof1Ctrl_19_oe = GEN_319;
  assign iof1Ctrl_19_ie = GEN_320;
  assign iof1Ctrl_20_oval = GEN_324;
  assign iof1Ctrl_20_oe = GEN_325;
  assign iof1Ctrl_20_ie = GEN_326;
  assign iof1Ctrl_21_oval = GEN_330;
  assign iof1Ctrl_21_oe = GEN_331;
  assign iof1Ctrl_21_ie = GEN_332;
  assign iof1Ctrl_22_oval = GEN_336;
  assign iof1Ctrl_22_oe = GEN_337;
  assign iof1Ctrl_22_ie = GEN_338;
  assign iof1Ctrl_23_oval = GEN_342;
  assign iof1Ctrl_23_oe = GEN_343;
  assign iof1Ctrl_23_ie = GEN_344;
  assign iof1Ctrl_24_oval = GEN_348;
  assign iof1Ctrl_24_oe = GEN_349;
  assign iof1Ctrl_24_ie = GEN_350;
  assign iof1Ctrl_25_oval = GEN_354;
  assign iof1Ctrl_25_oe = GEN_355;
  assign iof1Ctrl_25_ie = GEN_356;
  assign iof1Ctrl_26_oval = GEN_360;
  assign iof1Ctrl_26_oe = GEN_361;
  assign iof1Ctrl_26_ie = GEN_362;
  assign iof1Ctrl_27_oval = GEN_366;
  assign iof1Ctrl_27_oe = GEN_367;
  assign iof1Ctrl_27_ie = GEN_368;
  assign iof1Ctrl_28_oval = GEN_372;
  assign iof1Ctrl_28_oe = GEN_373;
  assign iof1Ctrl_28_ie = GEN_374;
  assign iof1Ctrl_29_oval = GEN_378;
  assign iof1Ctrl_29_oe = GEN_379;
  assign iof1Ctrl_29_ie = GEN_380;
  assign iof1Ctrl_30_oval = GEN_384;
  assign iof1Ctrl_30_oe = GEN_385;
  assign iof1Ctrl_30_ie = GEN_386;
  assign iof1Ctrl_31_oval = GEN_390;
  assign iof1Ctrl_31_oe = GEN_391;
  assign iof1Ctrl_31_ie = GEN_392;
  assign iofCtrl_0_oval = T_7575_oval;
  assign iofCtrl_0_oe = T_7575_oe;
  assign iofCtrl_0_ie = T_7575_ie;
  assign iofCtrl_1_oval = T_7611_oval;
  assign iofCtrl_1_oe = T_7611_oe;
  assign iofCtrl_1_ie = T_7611_ie;
  assign iofCtrl_2_oval = T_7647_oval;
  assign iofCtrl_2_oe = T_7647_oe;
  assign iofCtrl_2_ie = T_7647_ie;
  assign iofCtrl_3_oval = T_7683_oval;
  assign iofCtrl_3_oe = T_7683_oe;
  assign iofCtrl_3_ie = T_7683_ie;
  assign iofCtrl_4_oval = T_7719_oval;
  assign iofCtrl_4_oe = T_7719_oe;
  assign iofCtrl_4_ie = T_7719_ie;
  assign iofCtrl_5_oval = T_7755_oval;
  assign iofCtrl_5_oe = T_7755_oe;
  assign iofCtrl_5_ie = T_7755_ie;
  assign iofCtrl_6_oval = T_7791_oval;
  assign iofCtrl_6_oe = T_7791_oe;
  assign iofCtrl_6_ie = T_7791_ie;
  assign iofCtrl_7_oval = T_7827_oval;
  assign iofCtrl_7_oe = T_7827_oe;
  assign iofCtrl_7_ie = T_7827_ie;
  assign iofCtrl_8_oval = T_7863_oval;
  assign iofCtrl_8_oe = T_7863_oe;
  assign iofCtrl_8_ie = T_7863_ie;
  assign iofCtrl_9_oval = T_7899_oval;
  assign iofCtrl_9_oe = T_7899_oe;
  assign iofCtrl_9_ie = T_7899_ie;
  assign iofCtrl_10_oval = T_7935_oval;
  assign iofCtrl_10_oe = T_7935_oe;
  assign iofCtrl_10_ie = T_7935_ie;
  assign iofCtrl_11_oval = T_7971_oval;
  assign iofCtrl_11_oe = T_7971_oe;
  assign iofCtrl_11_ie = T_7971_ie;
  assign iofCtrl_12_oval = T_8007_oval;
  assign iofCtrl_12_oe = T_8007_oe;
  assign iofCtrl_12_ie = T_8007_ie;
  assign iofCtrl_13_oval = T_8043_oval;
  assign iofCtrl_13_oe = T_8043_oe;
  assign iofCtrl_13_ie = T_8043_ie;
  assign iofCtrl_14_oval = T_8079_oval;
  assign iofCtrl_14_oe = T_8079_oe;
  assign iofCtrl_14_ie = T_8079_ie;
  assign iofCtrl_15_oval = T_8115_oval;
  assign iofCtrl_15_oe = T_8115_oe;
  assign iofCtrl_15_ie = T_8115_ie;
  assign iofCtrl_16_oval = T_8151_oval;
  assign iofCtrl_16_oe = T_8151_oe;
  assign iofCtrl_16_ie = T_8151_ie;
  assign iofCtrl_17_oval = T_8187_oval;
  assign iofCtrl_17_oe = T_8187_oe;
  assign iofCtrl_17_ie = T_8187_ie;
  assign iofCtrl_18_oval = T_8223_oval;
  assign iofCtrl_18_oe = T_8223_oe;
  assign iofCtrl_18_ie = T_8223_ie;
  assign iofCtrl_19_oval = T_8259_oval;
  assign iofCtrl_19_oe = T_8259_oe;
  assign iofCtrl_19_ie = T_8259_ie;
  assign iofCtrl_20_oval = T_8295_oval;
  assign iofCtrl_20_oe = T_8295_oe;
  assign iofCtrl_20_ie = T_8295_ie;
  assign iofCtrl_21_oval = T_8331_oval;
  assign iofCtrl_21_oe = T_8331_oe;
  assign iofCtrl_21_ie = T_8331_ie;
  assign iofCtrl_22_oval = T_8367_oval;
  assign iofCtrl_22_oe = T_8367_oe;
  assign iofCtrl_22_ie = T_8367_ie;
  assign iofCtrl_23_oval = T_8403_oval;
  assign iofCtrl_23_oe = T_8403_oe;
  assign iofCtrl_23_ie = T_8403_ie;
  assign iofCtrl_24_oval = T_8439_oval;
  assign iofCtrl_24_oe = T_8439_oe;
  assign iofCtrl_24_ie = T_8439_ie;
  assign iofCtrl_25_oval = T_8475_oval;
  assign iofCtrl_25_oe = T_8475_oe;
  assign iofCtrl_25_ie = T_8475_ie;
  assign iofCtrl_26_oval = T_8511_oval;
  assign iofCtrl_26_oe = T_8511_oe;
  assign iofCtrl_26_ie = T_8511_ie;
  assign iofCtrl_27_oval = T_8547_oval;
  assign iofCtrl_27_oe = T_8547_oe;
  assign iofCtrl_27_ie = T_8547_ie;
  assign iofCtrl_28_oval = T_8583_oval;
  assign iofCtrl_28_oe = T_8583_oe;
  assign iofCtrl_28_ie = T_8583_ie;
  assign iofCtrl_29_oval = T_8619_oval;
  assign iofCtrl_29_oe = T_8619_oe;
  assign iofCtrl_29_ie = T_8619_ie;
  assign iofCtrl_30_oval = T_8655_oval;
  assign iofCtrl_30_oe = T_8655_oe;
  assign iofCtrl_30_ie = T_8655_ie;
  assign iofCtrl_31_oval = T_8691_oval;
  assign iofCtrl_31_oe = T_8691_oe;
  assign iofCtrl_31_ie = T_8691_ie;
  assign iofPlusSwPinCtrl_0_oval = iofCtrl_0_oval;
  assign iofPlusSwPinCtrl_0_oe = iofCtrl_0_oe;
  assign iofPlusSwPinCtrl_0_ie = iofCtrl_0_ie;
  assign iofPlusSwPinCtrl_0_pue = swPinCtrl_0_pue;
  assign iofPlusSwPinCtrl_0_ds = swPinCtrl_0_ds;
  assign iofPlusSwPinCtrl_1_oval = iofCtrl_1_oval;
  assign iofPlusSwPinCtrl_1_oe = iofCtrl_1_oe;
  assign iofPlusSwPinCtrl_1_ie = iofCtrl_1_ie;
  assign iofPlusSwPinCtrl_1_pue = swPinCtrl_1_pue;
  assign iofPlusSwPinCtrl_1_ds = swPinCtrl_1_ds;
  assign iofPlusSwPinCtrl_2_oval = iofCtrl_2_oval;
  assign iofPlusSwPinCtrl_2_oe = iofCtrl_2_oe;
  assign iofPlusSwPinCtrl_2_ie = iofCtrl_2_ie;
  assign iofPlusSwPinCtrl_2_pue = swPinCtrl_2_pue;
  assign iofPlusSwPinCtrl_2_ds = swPinCtrl_2_ds;
  assign iofPlusSwPinCtrl_3_oval = iofCtrl_3_oval;
  assign iofPlusSwPinCtrl_3_oe = iofCtrl_3_oe;
  assign iofPlusSwPinCtrl_3_ie = iofCtrl_3_ie;
  assign iofPlusSwPinCtrl_3_pue = swPinCtrl_3_pue;
  assign iofPlusSwPinCtrl_3_ds = swPinCtrl_3_ds;
  assign iofPlusSwPinCtrl_4_oval = iofCtrl_4_oval;
  assign iofPlusSwPinCtrl_4_oe = iofCtrl_4_oe;
  assign iofPlusSwPinCtrl_4_ie = iofCtrl_4_ie;
  assign iofPlusSwPinCtrl_4_pue = swPinCtrl_4_pue;
  assign iofPlusSwPinCtrl_4_ds = swPinCtrl_4_ds;
  assign iofPlusSwPinCtrl_5_oval = iofCtrl_5_oval;
  assign iofPlusSwPinCtrl_5_oe = iofCtrl_5_oe;
  assign iofPlusSwPinCtrl_5_ie = iofCtrl_5_ie;
  assign iofPlusSwPinCtrl_5_pue = swPinCtrl_5_pue;
  assign iofPlusSwPinCtrl_5_ds = swPinCtrl_5_ds;
  assign iofPlusSwPinCtrl_6_oval = iofCtrl_6_oval;
  assign iofPlusSwPinCtrl_6_oe = iofCtrl_6_oe;
  assign iofPlusSwPinCtrl_6_ie = iofCtrl_6_ie;
  assign iofPlusSwPinCtrl_6_pue = swPinCtrl_6_pue;
  assign iofPlusSwPinCtrl_6_ds = swPinCtrl_6_ds;
  assign iofPlusSwPinCtrl_7_oval = iofCtrl_7_oval;
  assign iofPlusSwPinCtrl_7_oe = iofCtrl_7_oe;
  assign iofPlusSwPinCtrl_7_ie = iofCtrl_7_ie;
  assign iofPlusSwPinCtrl_7_pue = swPinCtrl_7_pue;
  assign iofPlusSwPinCtrl_7_ds = swPinCtrl_7_ds;
  assign iofPlusSwPinCtrl_8_oval = iofCtrl_8_oval;
  assign iofPlusSwPinCtrl_8_oe = iofCtrl_8_oe;
  assign iofPlusSwPinCtrl_8_ie = iofCtrl_8_ie;
  assign iofPlusSwPinCtrl_8_pue = swPinCtrl_8_pue;
  assign iofPlusSwPinCtrl_8_ds = swPinCtrl_8_ds;
  assign iofPlusSwPinCtrl_9_oval = iofCtrl_9_oval;
  assign iofPlusSwPinCtrl_9_oe = iofCtrl_9_oe;
  assign iofPlusSwPinCtrl_9_ie = iofCtrl_9_ie;
  assign iofPlusSwPinCtrl_9_pue = swPinCtrl_9_pue;
  assign iofPlusSwPinCtrl_9_ds = swPinCtrl_9_ds;
  assign iofPlusSwPinCtrl_10_oval = iofCtrl_10_oval;
  assign iofPlusSwPinCtrl_10_oe = iofCtrl_10_oe;
  assign iofPlusSwPinCtrl_10_ie = iofCtrl_10_ie;
  assign iofPlusSwPinCtrl_10_pue = swPinCtrl_10_pue;
  assign iofPlusSwPinCtrl_10_ds = swPinCtrl_10_ds;
  assign iofPlusSwPinCtrl_11_oval = iofCtrl_11_oval;
  assign iofPlusSwPinCtrl_11_oe = iofCtrl_11_oe;
  assign iofPlusSwPinCtrl_11_ie = iofCtrl_11_ie;
  assign iofPlusSwPinCtrl_11_pue = swPinCtrl_11_pue;
  assign iofPlusSwPinCtrl_11_ds = swPinCtrl_11_ds;
  assign iofPlusSwPinCtrl_12_oval = iofCtrl_12_oval;
  assign iofPlusSwPinCtrl_12_oe = iofCtrl_12_oe;
  assign iofPlusSwPinCtrl_12_ie = iofCtrl_12_ie;
  assign iofPlusSwPinCtrl_12_pue = swPinCtrl_12_pue;
  assign iofPlusSwPinCtrl_12_ds = swPinCtrl_12_ds;
  assign iofPlusSwPinCtrl_13_oval = iofCtrl_13_oval;
  assign iofPlusSwPinCtrl_13_oe = iofCtrl_13_oe;
  assign iofPlusSwPinCtrl_13_ie = iofCtrl_13_ie;
  assign iofPlusSwPinCtrl_13_pue = swPinCtrl_13_pue;
  assign iofPlusSwPinCtrl_13_ds = swPinCtrl_13_ds;
  assign iofPlusSwPinCtrl_14_oval = iofCtrl_14_oval;
  assign iofPlusSwPinCtrl_14_oe = iofCtrl_14_oe;
  assign iofPlusSwPinCtrl_14_ie = iofCtrl_14_ie;
  assign iofPlusSwPinCtrl_14_pue = swPinCtrl_14_pue;
  assign iofPlusSwPinCtrl_14_ds = swPinCtrl_14_ds;
  assign iofPlusSwPinCtrl_15_oval = iofCtrl_15_oval;
  assign iofPlusSwPinCtrl_15_oe = iofCtrl_15_oe;
  assign iofPlusSwPinCtrl_15_ie = iofCtrl_15_ie;
  assign iofPlusSwPinCtrl_15_pue = swPinCtrl_15_pue;
  assign iofPlusSwPinCtrl_15_ds = swPinCtrl_15_ds;
  assign iofPlusSwPinCtrl_16_oval = iofCtrl_16_oval;
  assign iofPlusSwPinCtrl_16_oe = iofCtrl_16_oe;
  assign iofPlusSwPinCtrl_16_ie = iofCtrl_16_ie;
  assign iofPlusSwPinCtrl_16_pue = swPinCtrl_16_pue;
  assign iofPlusSwPinCtrl_16_ds = swPinCtrl_16_ds;
  assign iofPlusSwPinCtrl_17_oval = iofCtrl_17_oval;
  assign iofPlusSwPinCtrl_17_oe = iofCtrl_17_oe;
  assign iofPlusSwPinCtrl_17_ie = iofCtrl_17_ie;
  assign iofPlusSwPinCtrl_17_pue = swPinCtrl_17_pue;
  assign iofPlusSwPinCtrl_17_ds = swPinCtrl_17_ds;
  assign iofPlusSwPinCtrl_18_oval = iofCtrl_18_oval;
  assign iofPlusSwPinCtrl_18_oe = iofCtrl_18_oe;
  assign iofPlusSwPinCtrl_18_ie = iofCtrl_18_ie;
  assign iofPlusSwPinCtrl_18_pue = swPinCtrl_18_pue;
  assign iofPlusSwPinCtrl_18_ds = swPinCtrl_18_ds;
  assign iofPlusSwPinCtrl_19_oval = iofCtrl_19_oval;
  assign iofPlusSwPinCtrl_19_oe = iofCtrl_19_oe;
  assign iofPlusSwPinCtrl_19_ie = iofCtrl_19_ie;
  assign iofPlusSwPinCtrl_19_pue = swPinCtrl_19_pue;
  assign iofPlusSwPinCtrl_19_ds = swPinCtrl_19_ds;
  assign iofPlusSwPinCtrl_20_oval = iofCtrl_20_oval;
  assign iofPlusSwPinCtrl_20_oe = iofCtrl_20_oe;
  assign iofPlusSwPinCtrl_20_ie = iofCtrl_20_ie;
  assign iofPlusSwPinCtrl_20_pue = swPinCtrl_20_pue;
  assign iofPlusSwPinCtrl_20_ds = swPinCtrl_20_ds;
  assign iofPlusSwPinCtrl_21_oval = iofCtrl_21_oval;
  assign iofPlusSwPinCtrl_21_oe = iofCtrl_21_oe;
  assign iofPlusSwPinCtrl_21_ie = iofCtrl_21_ie;
  assign iofPlusSwPinCtrl_21_pue = swPinCtrl_21_pue;
  assign iofPlusSwPinCtrl_21_ds = swPinCtrl_21_ds;
  assign iofPlusSwPinCtrl_22_oval = iofCtrl_22_oval;
  assign iofPlusSwPinCtrl_22_oe = iofCtrl_22_oe;
  assign iofPlusSwPinCtrl_22_ie = iofCtrl_22_ie;
  assign iofPlusSwPinCtrl_22_pue = swPinCtrl_22_pue;
  assign iofPlusSwPinCtrl_22_ds = swPinCtrl_22_ds;
  assign iofPlusSwPinCtrl_23_oval = iofCtrl_23_oval;
  assign iofPlusSwPinCtrl_23_oe = iofCtrl_23_oe;
  assign iofPlusSwPinCtrl_23_ie = iofCtrl_23_ie;
  assign iofPlusSwPinCtrl_23_pue = swPinCtrl_23_pue;
  assign iofPlusSwPinCtrl_23_ds = swPinCtrl_23_ds;
  assign iofPlusSwPinCtrl_24_oval = iofCtrl_24_oval;
  assign iofPlusSwPinCtrl_24_oe = iofCtrl_24_oe;
  assign iofPlusSwPinCtrl_24_ie = iofCtrl_24_ie;
  assign iofPlusSwPinCtrl_24_pue = swPinCtrl_24_pue;
  assign iofPlusSwPinCtrl_24_ds = swPinCtrl_24_ds;
  assign iofPlusSwPinCtrl_25_oval = iofCtrl_25_oval;
  assign iofPlusSwPinCtrl_25_oe = iofCtrl_25_oe;
  assign iofPlusSwPinCtrl_25_ie = iofCtrl_25_ie;
  assign iofPlusSwPinCtrl_25_pue = swPinCtrl_25_pue;
  assign iofPlusSwPinCtrl_25_ds = swPinCtrl_25_ds;
  assign iofPlusSwPinCtrl_26_oval = iofCtrl_26_oval;
  assign iofPlusSwPinCtrl_26_oe = iofCtrl_26_oe;
  assign iofPlusSwPinCtrl_26_ie = iofCtrl_26_ie;
  assign iofPlusSwPinCtrl_26_pue = swPinCtrl_26_pue;
  assign iofPlusSwPinCtrl_26_ds = swPinCtrl_26_ds;
  assign iofPlusSwPinCtrl_27_oval = iofCtrl_27_oval;
  assign iofPlusSwPinCtrl_27_oe = iofCtrl_27_oe;
  assign iofPlusSwPinCtrl_27_ie = iofCtrl_27_ie;
  assign iofPlusSwPinCtrl_27_pue = swPinCtrl_27_pue;
  assign iofPlusSwPinCtrl_27_ds = swPinCtrl_27_ds;
  assign iofPlusSwPinCtrl_28_oval = iofCtrl_28_oval;
  assign iofPlusSwPinCtrl_28_oe = iofCtrl_28_oe;
  assign iofPlusSwPinCtrl_28_ie = iofCtrl_28_ie;
  assign iofPlusSwPinCtrl_28_pue = swPinCtrl_28_pue;
  assign iofPlusSwPinCtrl_28_ds = swPinCtrl_28_ds;
  assign iofPlusSwPinCtrl_29_oval = iofCtrl_29_oval;
  assign iofPlusSwPinCtrl_29_oe = iofCtrl_29_oe;
  assign iofPlusSwPinCtrl_29_ie = iofCtrl_29_ie;
  assign iofPlusSwPinCtrl_29_pue = swPinCtrl_29_pue;
  assign iofPlusSwPinCtrl_29_ds = swPinCtrl_29_ds;
  assign iofPlusSwPinCtrl_30_oval = iofCtrl_30_oval;
  assign iofPlusSwPinCtrl_30_oe = iofCtrl_30_oe;
  assign iofPlusSwPinCtrl_30_ie = iofCtrl_30_ie;
  assign iofPlusSwPinCtrl_30_pue = swPinCtrl_30_pue;
  assign iofPlusSwPinCtrl_30_ds = swPinCtrl_30_ds;
  assign iofPlusSwPinCtrl_31_oval = iofCtrl_31_oval;
  assign iofPlusSwPinCtrl_31_oe = iofCtrl_31_oe;
  assign iofPlusSwPinCtrl_31_ie = iofCtrl_31_ie;
  assign iofPlusSwPinCtrl_31_pue = swPinCtrl_31_pue;
  assign iofPlusSwPinCtrl_31_ds = swPinCtrl_31_ds;
  assign T_7569 = pueReg_io_q[0];
  assign T_7570 = portReg[0];
  assign T_7571 = oeReg_io_q[0];
  assign T_7572 = dsReg[0];
  assign T_7573 = ieReg_io_q[0];
  assign GEN_201 = io_port_iof_0_0_o_valid ? io_port_iof_0_0_o_oval : swPinCtrl_0_oval;
  assign GEN_202 = io_port_iof_0_0_o_valid ? io_port_iof_0_0_o_oe : swPinCtrl_0_oe;
  assign GEN_203 = io_port_iof_0_0_o_valid ? io_port_iof_0_0_o_ie : swPinCtrl_0_ie;
  assign GEN_204 = io_port_iof_1_0_o_valid ? io_port_iof_1_0_o_oval : swPinCtrl_0_oval;
  assign GEN_205 = io_port_iof_1_0_o_valid ? io_port_iof_1_0_o_oe : swPinCtrl_0_oe;
  assign GEN_206 = io_port_iof_1_0_o_valid ? io_port_iof_1_0_o_ie : swPinCtrl_0_ie;
  assign T_7574 = iofSelReg[0];
  assign T_7575_oval = T_7574 ? iof1Ctrl_0_oval : iof0Ctrl_0_oval;
  assign T_7575_oe = T_7574 ? iof1Ctrl_0_oe : iof0Ctrl_0_oe;
  assign T_7575_ie = T_7574 ? iof1Ctrl_0_ie : iof0Ctrl_0_ie;
  assign T_7579 = iofEnReg_io_q[0];
  assign T_7580_oval = T_7579 ? iofPlusSwPinCtrl_0_oval : swPinCtrl_0_oval;
  assign T_7580_oe = T_7579 ? iofPlusSwPinCtrl_0_oe : swPinCtrl_0_oe;
  assign T_7580_ie = T_7579 ? iofPlusSwPinCtrl_0_ie : swPinCtrl_0_ie;
  assign T_7580_pue = T_7579 ? iofPlusSwPinCtrl_0_pue : swPinCtrl_0_pue;
  assign T_7580_ds = T_7579 ? iofPlusSwPinCtrl_0_ds : swPinCtrl_0_ds;
  assign T_7586 = xorReg[0];
  assign T_7587 = T_7580_oval ^ T_7586;
  assign T_7588 = riseIpReg[0];
  assign T_7589 = riseIeReg[0];
  assign T_7590 = T_7588 & T_7589;
  assign T_7591 = fallIpReg[0];
  assign T_7592 = fallIeReg[0];
  assign T_7593 = T_7591 & T_7592;
  assign T_7594 = T_7590 | T_7593;
  assign T_7595 = highIpReg[0];
  assign T_7596 = highIeReg[0];
  assign T_7597 = T_7595 & T_7596;
  assign T_7598 = T_7594 | T_7597;
  assign T_7599 = lowIpReg[0];
  assign T_7600 = lowIeReg[0];
  assign T_7601 = T_7599 & T_7600;
  assign T_7602 = T_7598 | T_7601;
  assign T_7603 = inSyncReg[0];
  assign T_7605 = pueReg_io_q[1];
  assign T_7606 = portReg[1];
  assign T_7607 = oeReg_io_q[1];
  assign T_7608 = dsReg[1];
  assign T_7609 = ieReg_io_q[1];
  assign GEN_207 = io_port_iof_0_1_o_valid ? io_port_iof_0_1_o_oval : swPinCtrl_1_oval;
  assign GEN_208 = io_port_iof_0_1_o_valid ? io_port_iof_0_1_o_oe : swPinCtrl_1_oe;
  assign GEN_209 = io_port_iof_0_1_o_valid ? io_port_iof_0_1_o_ie : swPinCtrl_1_ie;
  assign GEN_210 = io_port_iof_1_1_o_valid ? io_port_iof_1_1_o_oval : swPinCtrl_1_oval;
  assign GEN_211 = io_port_iof_1_1_o_valid ? io_port_iof_1_1_o_oe : swPinCtrl_1_oe;
  assign GEN_212 = io_port_iof_1_1_o_valid ? io_port_iof_1_1_o_ie : swPinCtrl_1_ie;
  assign T_7610 = iofSelReg[1];
  assign T_7611_oval = T_7610 ? iof1Ctrl_1_oval : iof0Ctrl_1_oval;
  assign T_7611_oe = T_7610 ? iof1Ctrl_1_oe : iof0Ctrl_1_oe;
  assign T_7611_ie = T_7610 ? iof1Ctrl_1_ie : iof0Ctrl_1_ie;
  assign T_7615 = iofEnReg_io_q[1];
  assign T_7616_oval = T_7615 ? iofPlusSwPinCtrl_1_oval : swPinCtrl_1_oval;
  assign T_7616_oe = T_7615 ? iofPlusSwPinCtrl_1_oe : swPinCtrl_1_oe;
  assign T_7616_ie = T_7615 ? iofPlusSwPinCtrl_1_ie : swPinCtrl_1_ie;
  assign T_7616_pue = T_7615 ? iofPlusSwPinCtrl_1_pue : swPinCtrl_1_pue;
  assign T_7616_ds = T_7615 ? iofPlusSwPinCtrl_1_ds : swPinCtrl_1_ds;
  assign T_7622 = xorReg[1];
  assign T_7623 = T_7616_oval ^ T_7622;
  assign T_7624 = riseIpReg[1];
  assign T_7625 = riseIeReg[1];
  assign T_7626 = T_7624 & T_7625;
  assign T_7627 = fallIpReg[1];
  assign T_7628 = fallIeReg[1];
  assign T_7629 = T_7627 & T_7628;
  assign T_7630 = T_7626 | T_7629;
  assign T_7631 = highIpReg[1];
  assign T_7632 = highIeReg[1];
  assign T_7633 = T_7631 & T_7632;
  assign T_7634 = T_7630 | T_7633;
  assign T_7635 = lowIpReg[1];
  assign T_7636 = lowIeReg[1];
  assign T_7637 = T_7635 & T_7636;
  assign T_7638 = T_7634 | T_7637;
  assign T_7639 = inSyncReg[1];
  assign T_7641 = pueReg_io_q[2];
  assign T_7642 = portReg[2];
  assign T_7643 = oeReg_io_q[2];
  assign T_7644 = dsReg[2];
  assign T_7645 = ieReg_io_q[2];
  assign GEN_213 = io_port_iof_0_2_o_valid ? io_port_iof_0_2_o_oval : swPinCtrl_2_oval;
  assign GEN_214 = io_port_iof_0_2_o_valid ? io_port_iof_0_2_o_oe : swPinCtrl_2_oe;
  assign GEN_215 = io_port_iof_0_2_o_valid ? io_port_iof_0_2_o_ie : swPinCtrl_2_ie;
  assign GEN_216 = io_port_iof_1_2_o_valid ? io_port_iof_1_2_o_oval : swPinCtrl_2_oval;
  assign GEN_217 = io_port_iof_1_2_o_valid ? io_port_iof_1_2_o_oe : swPinCtrl_2_oe;
  assign GEN_218 = io_port_iof_1_2_o_valid ? io_port_iof_1_2_o_ie : swPinCtrl_2_ie;
  assign T_7646 = iofSelReg[2];
  assign T_7647_oval = T_7646 ? iof1Ctrl_2_oval : iof0Ctrl_2_oval;
  assign T_7647_oe = T_7646 ? iof1Ctrl_2_oe : iof0Ctrl_2_oe;
  assign T_7647_ie = T_7646 ? iof1Ctrl_2_ie : iof0Ctrl_2_ie;
  assign T_7651 = iofEnReg_io_q[2];
  assign T_7652_oval = T_7651 ? iofPlusSwPinCtrl_2_oval : swPinCtrl_2_oval;
  assign T_7652_oe = T_7651 ? iofPlusSwPinCtrl_2_oe : swPinCtrl_2_oe;
  assign T_7652_ie = T_7651 ? iofPlusSwPinCtrl_2_ie : swPinCtrl_2_ie;
  assign T_7652_pue = T_7651 ? iofPlusSwPinCtrl_2_pue : swPinCtrl_2_pue;
  assign T_7652_ds = T_7651 ? iofPlusSwPinCtrl_2_ds : swPinCtrl_2_ds;
  assign T_7658 = xorReg[2];
  assign T_7659 = T_7652_oval ^ T_7658;
  assign T_7660 = riseIpReg[2];
  assign T_7661 = riseIeReg[2];
  assign T_7662 = T_7660 & T_7661;
  assign T_7663 = fallIpReg[2];
  assign T_7664 = fallIeReg[2];
  assign T_7665 = T_7663 & T_7664;
  assign T_7666 = T_7662 | T_7665;
  assign T_7667 = highIpReg[2];
  assign T_7668 = highIeReg[2];
  assign T_7669 = T_7667 & T_7668;
  assign T_7670 = T_7666 | T_7669;
  assign T_7671 = lowIpReg[2];
  assign T_7672 = lowIeReg[2];
  assign T_7673 = T_7671 & T_7672;
  assign T_7674 = T_7670 | T_7673;
  assign T_7675 = inSyncReg[2];
  assign T_7677 = pueReg_io_q[3];
  assign T_7678 = portReg[3];
  assign T_7679 = oeReg_io_q[3];
  assign T_7680 = dsReg[3];
  assign T_7681 = ieReg_io_q[3];
  assign GEN_219 = io_port_iof_0_3_o_valid ? io_port_iof_0_3_o_oval : swPinCtrl_3_oval;
  assign GEN_220 = io_port_iof_0_3_o_valid ? io_port_iof_0_3_o_oe : swPinCtrl_3_oe;
  assign GEN_221 = io_port_iof_0_3_o_valid ? io_port_iof_0_3_o_ie : swPinCtrl_3_ie;
  assign GEN_222 = io_port_iof_1_3_o_valid ? io_port_iof_1_3_o_oval : swPinCtrl_3_oval;
  assign GEN_223 = io_port_iof_1_3_o_valid ? io_port_iof_1_3_o_oe : swPinCtrl_3_oe;
  assign GEN_224 = io_port_iof_1_3_o_valid ? io_port_iof_1_3_o_ie : swPinCtrl_3_ie;
  assign T_7682 = iofSelReg[3];
  assign T_7683_oval = T_7682 ? iof1Ctrl_3_oval : iof0Ctrl_3_oval;
  assign T_7683_oe = T_7682 ? iof1Ctrl_3_oe : iof0Ctrl_3_oe;
  assign T_7683_ie = T_7682 ? iof1Ctrl_3_ie : iof0Ctrl_3_ie;
  assign T_7687 = iofEnReg_io_q[3];
  assign T_7688_oval = T_7687 ? iofPlusSwPinCtrl_3_oval : swPinCtrl_3_oval;
  assign T_7688_oe = T_7687 ? iofPlusSwPinCtrl_3_oe : swPinCtrl_3_oe;
  assign T_7688_ie = T_7687 ? iofPlusSwPinCtrl_3_ie : swPinCtrl_3_ie;
  assign T_7688_pue = T_7687 ? iofPlusSwPinCtrl_3_pue : swPinCtrl_3_pue;
  assign T_7688_ds = T_7687 ? iofPlusSwPinCtrl_3_ds : swPinCtrl_3_ds;
  assign T_7694 = xorReg[3];
  assign T_7695 = T_7688_oval ^ T_7694;
  assign T_7696 = riseIpReg[3];
  assign T_7697 = riseIeReg[3];
  assign T_7698 = T_7696 & T_7697;
  assign T_7699 = fallIpReg[3];
  assign T_7700 = fallIeReg[3];
  assign T_7701 = T_7699 & T_7700;
  assign T_7702 = T_7698 | T_7701;
  assign T_7703 = highIpReg[3];
  assign T_7704 = highIeReg[3];
  assign T_7705 = T_7703 & T_7704;
  assign T_7706 = T_7702 | T_7705;
  assign T_7707 = lowIpReg[3];
  assign T_7708 = lowIeReg[3];
  assign T_7709 = T_7707 & T_7708;
  assign T_7710 = T_7706 | T_7709;
  assign T_7711 = inSyncReg[3];
  assign T_7713 = pueReg_io_q[4];
  assign T_7714 = portReg[4];
  assign T_7715 = oeReg_io_q[4];
  assign T_7716 = dsReg[4];
  assign T_7717 = ieReg_io_q[4];
  assign GEN_225 = io_port_iof_0_4_o_valid ? io_port_iof_0_4_o_oval : swPinCtrl_4_oval;
  assign GEN_226 = io_port_iof_0_4_o_valid ? io_port_iof_0_4_o_oe : swPinCtrl_4_oe;
  assign GEN_227 = io_port_iof_0_4_o_valid ? io_port_iof_0_4_o_ie : swPinCtrl_4_ie;
  assign GEN_228 = io_port_iof_1_4_o_valid ? io_port_iof_1_4_o_oval : swPinCtrl_4_oval;
  assign GEN_229 = io_port_iof_1_4_o_valid ? io_port_iof_1_4_o_oe : swPinCtrl_4_oe;
  assign GEN_230 = io_port_iof_1_4_o_valid ? io_port_iof_1_4_o_ie : swPinCtrl_4_ie;
  assign T_7718 = iofSelReg[4];
  assign T_7719_oval = T_7718 ? iof1Ctrl_4_oval : iof0Ctrl_4_oval;
  assign T_7719_oe = T_7718 ? iof1Ctrl_4_oe : iof0Ctrl_4_oe;
  assign T_7719_ie = T_7718 ? iof1Ctrl_4_ie : iof0Ctrl_4_ie;
  assign T_7723 = iofEnReg_io_q[4];
  assign T_7724_oval = T_7723 ? iofPlusSwPinCtrl_4_oval : swPinCtrl_4_oval;
  assign T_7724_oe = T_7723 ? iofPlusSwPinCtrl_4_oe : swPinCtrl_4_oe;
  assign T_7724_ie = T_7723 ? iofPlusSwPinCtrl_4_ie : swPinCtrl_4_ie;
  assign T_7724_pue = T_7723 ? iofPlusSwPinCtrl_4_pue : swPinCtrl_4_pue;
  assign T_7724_ds = T_7723 ? iofPlusSwPinCtrl_4_ds : swPinCtrl_4_ds;
  assign T_7730 = xorReg[4];
  assign T_7731 = T_7724_oval ^ T_7730;
  assign T_7732 = riseIpReg[4];
  assign T_7733 = riseIeReg[4];
  assign T_7734 = T_7732 & T_7733;
  assign T_7735 = fallIpReg[4];
  assign T_7736 = fallIeReg[4];
  assign T_7737 = T_7735 & T_7736;
  assign T_7738 = T_7734 | T_7737;
  assign T_7739 = highIpReg[4];
  assign T_7740 = highIeReg[4];
  assign T_7741 = T_7739 & T_7740;
  assign T_7742 = T_7738 | T_7741;
  assign T_7743 = lowIpReg[4];
  assign T_7744 = lowIeReg[4];
  assign T_7745 = T_7743 & T_7744;
  assign T_7746 = T_7742 | T_7745;
  assign T_7747 = inSyncReg[4];
  assign T_7749 = pueReg_io_q[5];
  assign T_7750 = portReg[5];
  assign T_7751 = oeReg_io_q[5];
  assign T_7752 = dsReg[5];
  assign T_7753 = ieReg_io_q[5];
  assign GEN_231 = io_port_iof_0_5_o_valid ? io_port_iof_0_5_o_oval : swPinCtrl_5_oval;
  assign GEN_232 = io_port_iof_0_5_o_valid ? io_port_iof_0_5_o_oe : swPinCtrl_5_oe;
  assign GEN_233 = io_port_iof_0_5_o_valid ? io_port_iof_0_5_o_ie : swPinCtrl_5_ie;
  assign GEN_234 = io_port_iof_1_5_o_valid ? io_port_iof_1_5_o_oval : swPinCtrl_5_oval;
  assign GEN_235 = io_port_iof_1_5_o_valid ? io_port_iof_1_5_o_oe : swPinCtrl_5_oe;
  assign GEN_236 = io_port_iof_1_5_o_valid ? io_port_iof_1_5_o_ie : swPinCtrl_5_ie;
  assign T_7754 = iofSelReg[5];
  assign T_7755_oval = T_7754 ? iof1Ctrl_5_oval : iof0Ctrl_5_oval;
  assign T_7755_oe = T_7754 ? iof1Ctrl_5_oe : iof0Ctrl_5_oe;
  assign T_7755_ie = T_7754 ? iof1Ctrl_5_ie : iof0Ctrl_5_ie;
  assign T_7759 = iofEnReg_io_q[5];
  assign T_7760_oval = T_7759 ? iofPlusSwPinCtrl_5_oval : swPinCtrl_5_oval;
  assign T_7760_oe = T_7759 ? iofPlusSwPinCtrl_5_oe : swPinCtrl_5_oe;
  assign T_7760_ie = T_7759 ? iofPlusSwPinCtrl_5_ie : swPinCtrl_5_ie;
  assign T_7760_pue = T_7759 ? iofPlusSwPinCtrl_5_pue : swPinCtrl_5_pue;
  assign T_7760_ds = T_7759 ? iofPlusSwPinCtrl_5_ds : swPinCtrl_5_ds;
  assign T_7766 = xorReg[5];
  assign T_7767 = T_7760_oval ^ T_7766;
  assign T_7768 = riseIpReg[5];
  assign T_7769 = riseIeReg[5];
  assign T_7770 = T_7768 & T_7769;
  assign T_7771 = fallIpReg[5];
  assign T_7772 = fallIeReg[5];
  assign T_7773 = T_7771 & T_7772;
  assign T_7774 = T_7770 | T_7773;
  assign T_7775 = highIpReg[5];
  assign T_7776 = highIeReg[5];
  assign T_7777 = T_7775 & T_7776;
  assign T_7778 = T_7774 | T_7777;
  assign T_7779 = lowIpReg[5];
  assign T_7780 = lowIeReg[5];
  assign T_7781 = T_7779 & T_7780;
  assign T_7782 = T_7778 | T_7781;
  assign T_7783 = inSyncReg[5];
  assign T_7785 = pueReg_io_q[6];
  assign T_7786 = portReg[6];
  assign T_7787 = oeReg_io_q[6];
  assign T_7788 = dsReg[6];
  assign T_7789 = ieReg_io_q[6];
  assign GEN_237 = io_port_iof_0_6_o_valid ? io_port_iof_0_6_o_oval : swPinCtrl_6_oval;
  assign GEN_238 = io_port_iof_0_6_o_valid ? io_port_iof_0_6_o_oe : swPinCtrl_6_oe;
  assign GEN_239 = io_port_iof_0_6_o_valid ? io_port_iof_0_6_o_ie : swPinCtrl_6_ie;
  assign GEN_240 = io_port_iof_1_6_o_valid ? io_port_iof_1_6_o_oval : swPinCtrl_6_oval;
  assign GEN_241 = io_port_iof_1_6_o_valid ? io_port_iof_1_6_o_oe : swPinCtrl_6_oe;
  assign GEN_242 = io_port_iof_1_6_o_valid ? io_port_iof_1_6_o_ie : swPinCtrl_6_ie;
  assign T_7790 = iofSelReg[6];
  assign T_7791_oval = T_7790 ? iof1Ctrl_6_oval : iof0Ctrl_6_oval;
  assign T_7791_oe = T_7790 ? iof1Ctrl_6_oe : iof0Ctrl_6_oe;
  assign T_7791_ie = T_7790 ? iof1Ctrl_6_ie : iof0Ctrl_6_ie;
  assign T_7795 = iofEnReg_io_q[6];
  assign T_7796_oval = T_7795 ? iofPlusSwPinCtrl_6_oval : swPinCtrl_6_oval;
  assign T_7796_oe = T_7795 ? iofPlusSwPinCtrl_6_oe : swPinCtrl_6_oe;
  assign T_7796_ie = T_7795 ? iofPlusSwPinCtrl_6_ie : swPinCtrl_6_ie;
  assign T_7796_pue = T_7795 ? iofPlusSwPinCtrl_6_pue : swPinCtrl_6_pue;
  assign T_7796_ds = T_7795 ? iofPlusSwPinCtrl_6_ds : swPinCtrl_6_ds;
  assign T_7802 = xorReg[6];
  assign T_7803 = T_7796_oval ^ T_7802;
  assign T_7804 = riseIpReg[6];
  assign T_7805 = riseIeReg[6];
  assign T_7806 = T_7804 & T_7805;
  assign T_7807 = fallIpReg[6];
  assign T_7808 = fallIeReg[6];
  assign T_7809 = T_7807 & T_7808;
  assign T_7810 = T_7806 | T_7809;
  assign T_7811 = highIpReg[6];
  assign T_7812 = highIeReg[6];
  assign T_7813 = T_7811 & T_7812;
  assign T_7814 = T_7810 | T_7813;
  assign T_7815 = lowIpReg[6];
  assign T_7816 = lowIeReg[6];
  assign T_7817 = T_7815 & T_7816;
  assign T_7818 = T_7814 | T_7817;
  assign T_7819 = inSyncReg[6];
  assign T_7821 = pueReg_io_q[7];
  assign T_7822 = portReg[7];
  assign T_7823 = oeReg_io_q[7];
  assign T_7824 = dsReg[7];
  assign T_7825 = ieReg_io_q[7];
  assign GEN_243 = io_port_iof_0_7_o_valid ? io_port_iof_0_7_o_oval : swPinCtrl_7_oval;
  assign GEN_244 = io_port_iof_0_7_o_valid ? io_port_iof_0_7_o_oe : swPinCtrl_7_oe;
  assign GEN_245 = io_port_iof_0_7_o_valid ? io_port_iof_0_7_o_ie : swPinCtrl_7_ie;
  assign GEN_246 = io_port_iof_1_7_o_valid ? io_port_iof_1_7_o_oval : swPinCtrl_7_oval;
  assign GEN_247 = io_port_iof_1_7_o_valid ? io_port_iof_1_7_o_oe : swPinCtrl_7_oe;
  assign GEN_248 = io_port_iof_1_7_o_valid ? io_port_iof_1_7_o_ie : swPinCtrl_7_ie;
  assign T_7826 = iofSelReg[7];
  assign T_7827_oval = T_7826 ? iof1Ctrl_7_oval : iof0Ctrl_7_oval;
  assign T_7827_oe = T_7826 ? iof1Ctrl_7_oe : iof0Ctrl_7_oe;
  assign T_7827_ie = T_7826 ? iof1Ctrl_7_ie : iof0Ctrl_7_ie;
  assign T_7831 = iofEnReg_io_q[7];
  assign T_7832_oval = T_7831 ? iofPlusSwPinCtrl_7_oval : swPinCtrl_7_oval;
  assign T_7832_oe = T_7831 ? iofPlusSwPinCtrl_7_oe : swPinCtrl_7_oe;
  assign T_7832_ie = T_7831 ? iofPlusSwPinCtrl_7_ie : swPinCtrl_7_ie;
  assign T_7832_pue = T_7831 ? iofPlusSwPinCtrl_7_pue : swPinCtrl_7_pue;
  assign T_7832_ds = T_7831 ? iofPlusSwPinCtrl_7_ds : swPinCtrl_7_ds;
  assign T_7838 = xorReg[7];
  assign T_7839 = T_7832_oval ^ T_7838;
  assign T_7840 = riseIpReg[7];
  assign T_7841 = riseIeReg[7];
  assign T_7842 = T_7840 & T_7841;
  assign T_7843 = fallIpReg[7];
  assign T_7844 = fallIeReg[7];
  assign T_7845 = T_7843 & T_7844;
  assign T_7846 = T_7842 | T_7845;
  assign T_7847 = highIpReg[7];
  assign T_7848 = highIeReg[7];
  assign T_7849 = T_7847 & T_7848;
  assign T_7850 = T_7846 | T_7849;
  assign T_7851 = lowIpReg[7];
  assign T_7852 = lowIeReg[7];
  assign T_7853 = T_7851 & T_7852;
  assign T_7854 = T_7850 | T_7853;
  assign T_7855 = inSyncReg[7];
  assign T_7857 = pueReg_io_q[8];
  assign T_7858 = portReg[8];
  assign T_7859 = oeReg_io_q[8];
  assign T_7860 = dsReg[8];
  assign T_7861 = ieReg_io_q[8];
  assign GEN_249 = io_port_iof_0_8_o_valid ? io_port_iof_0_8_o_oval : swPinCtrl_8_oval;
  assign GEN_250 = io_port_iof_0_8_o_valid ? io_port_iof_0_8_o_oe : swPinCtrl_8_oe;
  assign GEN_251 = io_port_iof_0_8_o_valid ? io_port_iof_0_8_o_ie : swPinCtrl_8_ie;
  assign GEN_252 = io_port_iof_1_8_o_valid ? io_port_iof_1_8_o_oval : swPinCtrl_8_oval;
  assign GEN_253 = io_port_iof_1_8_o_valid ? io_port_iof_1_8_o_oe : swPinCtrl_8_oe;
  assign GEN_254 = io_port_iof_1_8_o_valid ? io_port_iof_1_8_o_ie : swPinCtrl_8_ie;
  assign T_7862 = iofSelReg[8];
  assign T_7863_oval = T_7862 ? iof1Ctrl_8_oval : iof0Ctrl_8_oval;
  assign T_7863_oe = T_7862 ? iof1Ctrl_8_oe : iof0Ctrl_8_oe;
  assign T_7863_ie = T_7862 ? iof1Ctrl_8_ie : iof0Ctrl_8_ie;
  assign T_7867 = iofEnReg_io_q[8];
  assign T_7868_oval = T_7867 ? iofPlusSwPinCtrl_8_oval : swPinCtrl_8_oval;
  assign T_7868_oe = T_7867 ? iofPlusSwPinCtrl_8_oe : swPinCtrl_8_oe;
  assign T_7868_ie = T_7867 ? iofPlusSwPinCtrl_8_ie : swPinCtrl_8_ie;
  assign T_7868_pue = T_7867 ? iofPlusSwPinCtrl_8_pue : swPinCtrl_8_pue;
  assign T_7868_ds = T_7867 ? iofPlusSwPinCtrl_8_ds : swPinCtrl_8_ds;
  assign T_7874 = xorReg[8];
  assign T_7875 = T_7868_oval ^ T_7874;
  assign T_7876 = riseIpReg[8];
  assign T_7877 = riseIeReg[8];
  assign T_7878 = T_7876 & T_7877;
  assign T_7879 = fallIpReg[8];
  assign T_7880 = fallIeReg[8];
  assign T_7881 = T_7879 & T_7880;
  assign T_7882 = T_7878 | T_7881;
  assign T_7883 = highIpReg[8];
  assign T_7884 = highIeReg[8];
  assign T_7885 = T_7883 & T_7884;
  assign T_7886 = T_7882 | T_7885;
  assign T_7887 = lowIpReg[8];
  assign T_7888 = lowIeReg[8];
  assign T_7889 = T_7887 & T_7888;
  assign T_7890 = T_7886 | T_7889;
  assign T_7891 = inSyncReg[8];
  assign T_7893 = pueReg_io_q[9];
  assign T_7894 = portReg[9];
  assign T_7895 = oeReg_io_q[9];
  assign T_7896 = dsReg[9];
  assign T_7897 = ieReg_io_q[9];
  assign GEN_255 = io_port_iof_0_9_o_valid ? io_port_iof_0_9_o_oval : swPinCtrl_9_oval;
  assign GEN_256 = io_port_iof_0_9_o_valid ? io_port_iof_0_9_o_oe : swPinCtrl_9_oe;
  assign GEN_257 = io_port_iof_0_9_o_valid ? io_port_iof_0_9_o_ie : swPinCtrl_9_ie;
  assign GEN_258 = io_port_iof_1_9_o_valid ? io_port_iof_1_9_o_oval : swPinCtrl_9_oval;
  assign GEN_259 = io_port_iof_1_9_o_valid ? io_port_iof_1_9_o_oe : swPinCtrl_9_oe;
  assign GEN_260 = io_port_iof_1_9_o_valid ? io_port_iof_1_9_o_ie : swPinCtrl_9_ie;
  assign T_7898 = iofSelReg[9];
  assign T_7899_oval = T_7898 ? iof1Ctrl_9_oval : iof0Ctrl_9_oval;
  assign T_7899_oe = T_7898 ? iof1Ctrl_9_oe : iof0Ctrl_9_oe;
  assign T_7899_ie = T_7898 ? iof1Ctrl_9_ie : iof0Ctrl_9_ie;
  assign T_7903 = iofEnReg_io_q[9];
  assign T_7904_oval = T_7903 ? iofPlusSwPinCtrl_9_oval : swPinCtrl_9_oval;
  assign T_7904_oe = T_7903 ? iofPlusSwPinCtrl_9_oe : swPinCtrl_9_oe;
  assign T_7904_ie = T_7903 ? iofPlusSwPinCtrl_9_ie : swPinCtrl_9_ie;
  assign T_7904_pue = T_7903 ? iofPlusSwPinCtrl_9_pue : swPinCtrl_9_pue;
  assign T_7904_ds = T_7903 ? iofPlusSwPinCtrl_9_ds : swPinCtrl_9_ds;
  assign T_7910 = xorReg[9];
  assign T_7911 = T_7904_oval ^ T_7910;
  assign T_7912 = riseIpReg[9];
  assign T_7913 = riseIeReg[9];
  assign T_7914 = T_7912 & T_7913;
  assign T_7915 = fallIpReg[9];
  assign T_7916 = fallIeReg[9];
  assign T_7917 = T_7915 & T_7916;
  assign T_7918 = T_7914 | T_7917;
  assign T_7919 = highIpReg[9];
  assign T_7920 = highIeReg[9];
  assign T_7921 = T_7919 & T_7920;
  assign T_7922 = T_7918 | T_7921;
  assign T_7923 = lowIpReg[9];
  assign T_7924 = lowIeReg[9];
  assign T_7925 = T_7923 & T_7924;
  assign T_7926 = T_7922 | T_7925;
  assign T_7927 = inSyncReg[9];
  assign T_7929 = pueReg_io_q[10];
  assign T_7930 = portReg[10];
  assign T_7931 = oeReg_io_q[10];
  assign T_7932 = dsReg[10];
  assign T_7933 = ieReg_io_q[10];
  assign GEN_261 = io_port_iof_0_10_o_valid ? io_port_iof_0_10_o_oval : swPinCtrl_10_oval;
  assign GEN_262 = io_port_iof_0_10_o_valid ? io_port_iof_0_10_o_oe : swPinCtrl_10_oe;
  assign GEN_263 = io_port_iof_0_10_o_valid ? io_port_iof_0_10_o_ie : swPinCtrl_10_ie;
  assign GEN_264 = io_port_iof_1_10_o_valid ? io_port_iof_1_10_o_oval : swPinCtrl_10_oval;
  assign GEN_265 = io_port_iof_1_10_o_valid ? io_port_iof_1_10_o_oe : swPinCtrl_10_oe;
  assign GEN_266 = io_port_iof_1_10_o_valid ? io_port_iof_1_10_o_ie : swPinCtrl_10_ie;
  assign T_7934 = iofSelReg[10];
  assign T_7935_oval = T_7934 ? iof1Ctrl_10_oval : iof0Ctrl_10_oval;
  assign T_7935_oe = T_7934 ? iof1Ctrl_10_oe : iof0Ctrl_10_oe;
  assign T_7935_ie = T_7934 ? iof1Ctrl_10_ie : iof0Ctrl_10_ie;
  assign T_7939 = iofEnReg_io_q[10];
  assign T_7940_oval = T_7939 ? iofPlusSwPinCtrl_10_oval : swPinCtrl_10_oval;
  assign T_7940_oe = T_7939 ? iofPlusSwPinCtrl_10_oe : swPinCtrl_10_oe;
  assign T_7940_ie = T_7939 ? iofPlusSwPinCtrl_10_ie : swPinCtrl_10_ie;
  assign T_7940_pue = T_7939 ? iofPlusSwPinCtrl_10_pue : swPinCtrl_10_pue;
  assign T_7940_ds = T_7939 ? iofPlusSwPinCtrl_10_ds : swPinCtrl_10_ds;
  assign T_7946 = xorReg[10];
  assign T_7947 = T_7940_oval ^ T_7946;
  assign T_7948 = riseIpReg[10];
  assign T_7949 = riseIeReg[10];
  assign T_7950 = T_7948 & T_7949;
  assign T_7951 = fallIpReg[10];
  assign T_7952 = fallIeReg[10];
  assign T_7953 = T_7951 & T_7952;
  assign T_7954 = T_7950 | T_7953;
  assign T_7955 = highIpReg[10];
  assign T_7956 = highIeReg[10];
  assign T_7957 = T_7955 & T_7956;
  assign T_7958 = T_7954 | T_7957;
  assign T_7959 = lowIpReg[10];
  assign T_7960 = lowIeReg[10];
  assign T_7961 = T_7959 & T_7960;
  assign T_7962 = T_7958 | T_7961;
  assign T_7963 = inSyncReg[10];
  assign T_7965 = pueReg_io_q[11];
  assign T_7966 = portReg[11];
  assign T_7967 = oeReg_io_q[11];
  assign T_7968 = dsReg[11];
  assign T_7969 = ieReg_io_q[11];
  assign GEN_267 = io_port_iof_0_11_o_valid ? io_port_iof_0_11_o_oval : swPinCtrl_11_oval;
  assign GEN_268 = io_port_iof_0_11_o_valid ? io_port_iof_0_11_o_oe : swPinCtrl_11_oe;
  assign GEN_269 = io_port_iof_0_11_o_valid ? io_port_iof_0_11_o_ie : swPinCtrl_11_ie;
  assign GEN_270 = io_port_iof_1_11_o_valid ? io_port_iof_1_11_o_oval : swPinCtrl_11_oval;
  assign GEN_271 = io_port_iof_1_11_o_valid ? io_port_iof_1_11_o_oe : swPinCtrl_11_oe;
  assign GEN_272 = io_port_iof_1_11_o_valid ? io_port_iof_1_11_o_ie : swPinCtrl_11_ie;
  assign T_7970 = iofSelReg[11];
  assign T_7971_oval = T_7970 ? iof1Ctrl_11_oval : iof0Ctrl_11_oval;
  assign T_7971_oe = T_7970 ? iof1Ctrl_11_oe : iof0Ctrl_11_oe;
  assign T_7971_ie = T_7970 ? iof1Ctrl_11_ie : iof0Ctrl_11_ie;
  assign T_7975 = iofEnReg_io_q[11];
  assign T_7976_oval = T_7975 ? iofPlusSwPinCtrl_11_oval : swPinCtrl_11_oval;
  assign T_7976_oe = T_7975 ? iofPlusSwPinCtrl_11_oe : swPinCtrl_11_oe;
  assign T_7976_ie = T_7975 ? iofPlusSwPinCtrl_11_ie : swPinCtrl_11_ie;
  assign T_7976_pue = T_7975 ? iofPlusSwPinCtrl_11_pue : swPinCtrl_11_pue;
  assign T_7976_ds = T_7975 ? iofPlusSwPinCtrl_11_ds : swPinCtrl_11_ds;
  assign T_7982 = xorReg[11];
  assign T_7983 = T_7976_oval ^ T_7982;
  assign T_7984 = riseIpReg[11];
  assign T_7985 = riseIeReg[11];
  assign T_7986 = T_7984 & T_7985;
  assign T_7987 = fallIpReg[11];
  assign T_7988 = fallIeReg[11];
  assign T_7989 = T_7987 & T_7988;
  assign T_7990 = T_7986 | T_7989;
  assign T_7991 = highIpReg[11];
  assign T_7992 = highIeReg[11];
  assign T_7993 = T_7991 & T_7992;
  assign T_7994 = T_7990 | T_7993;
  assign T_7995 = lowIpReg[11];
  assign T_7996 = lowIeReg[11];
  assign T_7997 = T_7995 & T_7996;
  assign T_7998 = T_7994 | T_7997;
  assign T_7999 = inSyncReg[11];
  assign T_8001 = pueReg_io_q[12];
  assign T_8002 = portReg[12];
  assign T_8003 = oeReg_io_q[12];
  assign T_8004 = dsReg[12];
  assign T_8005 = ieReg_io_q[12];
  assign GEN_273 = io_port_iof_0_12_o_valid ? io_port_iof_0_12_o_oval : swPinCtrl_12_oval;
  assign GEN_274 = io_port_iof_0_12_o_valid ? io_port_iof_0_12_o_oe : swPinCtrl_12_oe;
  assign GEN_275 = io_port_iof_0_12_o_valid ? io_port_iof_0_12_o_ie : swPinCtrl_12_ie;
  assign GEN_276 = io_port_iof_1_12_o_valid ? io_port_iof_1_12_o_oval : swPinCtrl_12_oval;
  assign GEN_277 = io_port_iof_1_12_o_valid ? io_port_iof_1_12_o_oe : swPinCtrl_12_oe;
  assign GEN_278 = io_port_iof_1_12_o_valid ? io_port_iof_1_12_o_ie : swPinCtrl_12_ie;
  assign T_8006 = iofSelReg[12];
  assign T_8007_oval = T_8006 ? iof1Ctrl_12_oval : iof0Ctrl_12_oval;
  assign T_8007_oe = T_8006 ? iof1Ctrl_12_oe : iof0Ctrl_12_oe;
  assign T_8007_ie = T_8006 ? iof1Ctrl_12_ie : iof0Ctrl_12_ie;
  assign T_8011 = iofEnReg_io_q[12];
  assign T_8012_oval = T_8011 ? iofPlusSwPinCtrl_12_oval : swPinCtrl_12_oval;
  assign T_8012_oe = T_8011 ? iofPlusSwPinCtrl_12_oe : swPinCtrl_12_oe;
  assign T_8012_ie = T_8011 ? iofPlusSwPinCtrl_12_ie : swPinCtrl_12_ie;
  assign T_8012_pue = T_8011 ? iofPlusSwPinCtrl_12_pue : swPinCtrl_12_pue;
  assign T_8012_ds = T_8011 ? iofPlusSwPinCtrl_12_ds : swPinCtrl_12_ds;
  assign T_8018 = xorReg[12];
  assign T_8019 = T_8012_oval ^ T_8018;
  assign T_8020 = riseIpReg[12];
  assign T_8021 = riseIeReg[12];
  assign T_8022 = T_8020 & T_8021;
  assign T_8023 = fallIpReg[12];
  assign T_8024 = fallIeReg[12];
  assign T_8025 = T_8023 & T_8024;
  assign T_8026 = T_8022 | T_8025;
  assign T_8027 = highIpReg[12];
  assign T_8028 = highIeReg[12];
  assign T_8029 = T_8027 & T_8028;
  assign T_8030 = T_8026 | T_8029;
  assign T_8031 = lowIpReg[12];
  assign T_8032 = lowIeReg[12];
  assign T_8033 = T_8031 & T_8032;
  assign T_8034 = T_8030 | T_8033;
  assign T_8035 = inSyncReg[12];
  assign T_8037 = pueReg_io_q[13];
  assign T_8038 = portReg[13];
  assign T_8039 = oeReg_io_q[13];
  assign T_8040 = dsReg[13];
  assign T_8041 = ieReg_io_q[13];
  assign GEN_279 = io_port_iof_0_13_o_valid ? io_port_iof_0_13_o_oval : swPinCtrl_13_oval;
  assign GEN_280 = io_port_iof_0_13_o_valid ? io_port_iof_0_13_o_oe : swPinCtrl_13_oe;
  assign GEN_281 = io_port_iof_0_13_o_valid ? io_port_iof_0_13_o_ie : swPinCtrl_13_ie;
  assign GEN_282 = io_port_iof_1_13_o_valid ? io_port_iof_1_13_o_oval : swPinCtrl_13_oval;
  assign GEN_283 = io_port_iof_1_13_o_valid ? io_port_iof_1_13_o_oe : swPinCtrl_13_oe;
  assign GEN_284 = io_port_iof_1_13_o_valid ? io_port_iof_1_13_o_ie : swPinCtrl_13_ie;
  assign T_8042 = iofSelReg[13];
  assign T_8043_oval = T_8042 ? iof1Ctrl_13_oval : iof0Ctrl_13_oval;
  assign T_8043_oe = T_8042 ? iof1Ctrl_13_oe : iof0Ctrl_13_oe;
  assign T_8043_ie = T_8042 ? iof1Ctrl_13_ie : iof0Ctrl_13_ie;
  assign T_8047 = iofEnReg_io_q[13];
  assign T_8048_oval = T_8047 ? iofPlusSwPinCtrl_13_oval : swPinCtrl_13_oval;
  assign T_8048_oe = T_8047 ? iofPlusSwPinCtrl_13_oe : swPinCtrl_13_oe;
  assign T_8048_ie = T_8047 ? iofPlusSwPinCtrl_13_ie : swPinCtrl_13_ie;
  assign T_8048_pue = T_8047 ? iofPlusSwPinCtrl_13_pue : swPinCtrl_13_pue;
  assign T_8048_ds = T_8047 ? iofPlusSwPinCtrl_13_ds : swPinCtrl_13_ds;
  assign T_8054 = xorReg[13];
  assign T_8055 = T_8048_oval ^ T_8054;
  assign T_8056 = riseIpReg[13];
  assign T_8057 = riseIeReg[13];
  assign T_8058 = T_8056 & T_8057;
  assign T_8059 = fallIpReg[13];
  assign T_8060 = fallIeReg[13];
  assign T_8061 = T_8059 & T_8060;
  assign T_8062 = T_8058 | T_8061;
  assign T_8063 = highIpReg[13];
  assign T_8064 = highIeReg[13];
  assign T_8065 = T_8063 & T_8064;
  assign T_8066 = T_8062 | T_8065;
  assign T_8067 = lowIpReg[13];
  assign T_8068 = lowIeReg[13];
  assign T_8069 = T_8067 & T_8068;
  assign T_8070 = T_8066 | T_8069;
  assign T_8071 = inSyncReg[13];
  assign T_8073 = pueReg_io_q[14];
  assign T_8074 = portReg[14];
  assign T_8075 = oeReg_io_q[14];
  assign T_8076 = dsReg[14];
  assign T_8077 = ieReg_io_q[14];
  assign GEN_285 = io_port_iof_0_14_o_valid ? io_port_iof_0_14_o_oval : swPinCtrl_14_oval;
  assign GEN_286 = io_port_iof_0_14_o_valid ? io_port_iof_0_14_o_oe : swPinCtrl_14_oe;
  assign GEN_287 = io_port_iof_0_14_o_valid ? io_port_iof_0_14_o_ie : swPinCtrl_14_ie;
  assign GEN_288 = io_port_iof_1_14_o_valid ? io_port_iof_1_14_o_oval : swPinCtrl_14_oval;
  assign GEN_289 = io_port_iof_1_14_o_valid ? io_port_iof_1_14_o_oe : swPinCtrl_14_oe;
  assign GEN_290 = io_port_iof_1_14_o_valid ? io_port_iof_1_14_o_ie : swPinCtrl_14_ie;
  assign T_8078 = iofSelReg[14];
  assign T_8079_oval = T_8078 ? iof1Ctrl_14_oval : iof0Ctrl_14_oval;
  assign T_8079_oe = T_8078 ? iof1Ctrl_14_oe : iof0Ctrl_14_oe;
  assign T_8079_ie = T_8078 ? iof1Ctrl_14_ie : iof0Ctrl_14_ie;
  assign T_8083 = iofEnReg_io_q[14];
  assign T_8084_oval = T_8083 ? iofPlusSwPinCtrl_14_oval : swPinCtrl_14_oval;
  assign T_8084_oe = T_8083 ? iofPlusSwPinCtrl_14_oe : swPinCtrl_14_oe;
  assign T_8084_ie = T_8083 ? iofPlusSwPinCtrl_14_ie : swPinCtrl_14_ie;
  assign T_8084_pue = T_8083 ? iofPlusSwPinCtrl_14_pue : swPinCtrl_14_pue;
  assign T_8084_ds = T_8083 ? iofPlusSwPinCtrl_14_ds : swPinCtrl_14_ds;
  assign T_8090 = xorReg[14];
  assign T_8091 = T_8084_oval ^ T_8090;
  assign T_8092 = riseIpReg[14];
  assign T_8093 = riseIeReg[14];
  assign T_8094 = T_8092 & T_8093;
  assign T_8095 = fallIpReg[14];
  assign T_8096 = fallIeReg[14];
  assign T_8097 = T_8095 & T_8096;
  assign T_8098 = T_8094 | T_8097;
  assign T_8099 = highIpReg[14];
  assign T_8100 = highIeReg[14];
  assign T_8101 = T_8099 & T_8100;
  assign T_8102 = T_8098 | T_8101;
  assign T_8103 = lowIpReg[14];
  assign T_8104 = lowIeReg[14];
  assign T_8105 = T_8103 & T_8104;
  assign T_8106 = T_8102 | T_8105;
  assign T_8107 = inSyncReg[14];
  assign T_8109 = pueReg_io_q[15];
  assign T_8110 = portReg[15];
  assign T_8111 = oeReg_io_q[15];
  assign T_8112 = dsReg[15];
  assign T_8113 = ieReg_io_q[15];
  assign GEN_291 = io_port_iof_0_15_o_valid ? io_port_iof_0_15_o_oval : swPinCtrl_15_oval;
  assign GEN_292 = io_port_iof_0_15_o_valid ? io_port_iof_0_15_o_oe : swPinCtrl_15_oe;
  assign GEN_293 = io_port_iof_0_15_o_valid ? io_port_iof_0_15_o_ie : swPinCtrl_15_ie;
  assign GEN_294 = io_port_iof_1_15_o_valid ? io_port_iof_1_15_o_oval : swPinCtrl_15_oval;
  assign GEN_295 = io_port_iof_1_15_o_valid ? io_port_iof_1_15_o_oe : swPinCtrl_15_oe;
  assign GEN_296 = io_port_iof_1_15_o_valid ? io_port_iof_1_15_o_ie : swPinCtrl_15_ie;
  assign T_8114 = iofSelReg[15];
  assign T_8115_oval = T_8114 ? iof1Ctrl_15_oval : iof0Ctrl_15_oval;
  assign T_8115_oe = T_8114 ? iof1Ctrl_15_oe : iof0Ctrl_15_oe;
  assign T_8115_ie = T_8114 ? iof1Ctrl_15_ie : iof0Ctrl_15_ie;
  assign T_8119 = iofEnReg_io_q[15];
  assign T_8120_oval = T_8119 ? iofPlusSwPinCtrl_15_oval : swPinCtrl_15_oval;
  assign T_8120_oe = T_8119 ? iofPlusSwPinCtrl_15_oe : swPinCtrl_15_oe;
  assign T_8120_ie = T_8119 ? iofPlusSwPinCtrl_15_ie : swPinCtrl_15_ie;
  assign T_8120_pue = T_8119 ? iofPlusSwPinCtrl_15_pue : swPinCtrl_15_pue;
  assign T_8120_ds = T_8119 ? iofPlusSwPinCtrl_15_ds : swPinCtrl_15_ds;
  assign T_8126 = xorReg[15];
  assign T_8127 = T_8120_oval ^ T_8126;
  assign T_8128 = riseIpReg[15];
  assign T_8129 = riseIeReg[15];
  assign T_8130 = T_8128 & T_8129;
  assign T_8131 = fallIpReg[15];
  assign T_8132 = fallIeReg[15];
  assign T_8133 = T_8131 & T_8132;
  assign T_8134 = T_8130 | T_8133;
  assign T_8135 = highIpReg[15];
  assign T_8136 = highIeReg[15];
  assign T_8137 = T_8135 & T_8136;
  assign T_8138 = T_8134 | T_8137;
  assign T_8139 = lowIpReg[15];
  assign T_8140 = lowIeReg[15];
  assign T_8141 = T_8139 & T_8140;
  assign T_8142 = T_8138 | T_8141;
  assign T_8143 = inSyncReg[15];
  assign T_8145 = pueReg_io_q[16];
  assign T_8146 = portReg[16];
  assign T_8147 = oeReg_io_q[16];
  assign T_8148 = dsReg[16];
  assign T_8149 = ieReg_io_q[16];
  assign GEN_297 = io_port_iof_0_16_o_valid ? io_port_iof_0_16_o_oval : swPinCtrl_16_oval;
  assign GEN_298 = io_port_iof_0_16_o_valid ? io_port_iof_0_16_o_oe : swPinCtrl_16_oe;
  assign GEN_299 = io_port_iof_0_16_o_valid ? io_port_iof_0_16_o_ie : swPinCtrl_16_ie;
  assign GEN_300 = io_port_iof_1_16_o_valid ? io_port_iof_1_16_o_oval : swPinCtrl_16_oval;
  assign GEN_301 = io_port_iof_1_16_o_valid ? io_port_iof_1_16_o_oe : swPinCtrl_16_oe;
  assign GEN_302 = io_port_iof_1_16_o_valid ? io_port_iof_1_16_o_ie : swPinCtrl_16_ie;
  assign T_8150 = iofSelReg[16];
  assign T_8151_oval = T_8150 ? iof1Ctrl_16_oval : iof0Ctrl_16_oval;
  assign T_8151_oe = T_8150 ? iof1Ctrl_16_oe : iof0Ctrl_16_oe;
  assign T_8151_ie = T_8150 ? iof1Ctrl_16_ie : iof0Ctrl_16_ie;
  assign T_8155 = iofEnReg_io_q[16];
  assign T_8156_oval = T_8155 ? iofPlusSwPinCtrl_16_oval : swPinCtrl_16_oval;
  assign T_8156_oe = T_8155 ? iofPlusSwPinCtrl_16_oe : swPinCtrl_16_oe;
  assign T_8156_ie = T_8155 ? iofPlusSwPinCtrl_16_ie : swPinCtrl_16_ie;
  assign T_8156_pue = T_8155 ? iofPlusSwPinCtrl_16_pue : swPinCtrl_16_pue;
  assign T_8156_ds = T_8155 ? iofPlusSwPinCtrl_16_ds : swPinCtrl_16_ds;
  assign T_8162 = xorReg[16];
  assign T_8163 = T_8156_oval ^ T_8162;
  assign T_8164 = riseIpReg[16];
  assign T_8165 = riseIeReg[16];
  assign T_8166 = T_8164 & T_8165;
  assign T_8167 = fallIpReg[16];
  assign T_8168 = fallIeReg[16];
  assign T_8169 = T_8167 & T_8168;
  assign T_8170 = T_8166 | T_8169;
  assign T_8171 = highIpReg[16];
  assign T_8172 = highIeReg[16];
  assign T_8173 = T_8171 & T_8172;
  assign T_8174 = T_8170 | T_8173;
  assign T_8175 = lowIpReg[16];
  assign T_8176 = lowIeReg[16];
  assign T_8177 = T_8175 & T_8176;
  assign T_8178 = T_8174 | T_8177;
  assign T_8179 = inSyncReg[16];
  assign T_8181 = pueReg_io_q[17];
  assign T_8182 = portReg[17];
  assign T_8183 = oeReg_io_q[17];
  assign T_8184 = dsReg[17];
  assign T_8185 = ieReg_io_q[17];
  assign GEN_303 = io_port_iof_0_17_o_valid ? io_port_iof_0_17_o_oval : swPinCtrl_17_oval;
  assign GEN_304 = io_port_iof_0_17_o_valid ? io_port_iof_0_17_o_oe : swPinCtrl_17_oe;
  assign GEN_305 = io_port_iof_0_17_o_valid ? io_port_iof_0_17_o_ie : swPinCtrl_17_ie;
  assign GEN_306 = io_port_iof_1_17_o_valid ? io_port_iof_1_17_o_oval : swPinCtrl_17_oval;
  assign GEN_307 = io_port_iof_1_17_o_valid ? io_port_iof_1_17_o_oe : swPinCtrl_17_oe;
  assign GEN_308 = io_port_iof_1_17_o_valid ? io_port_iof_1_17_o_ie : swPinCtrl_17_ie;
  assign T_8186 = iofSelReg[17];
  assign T_8187_oval = T_8186 ? iof1Ctrl_17_oval : iof0Ctrl_17_oval;
  assign T_8187_oe = T_8186 ? iof1Ctrl_17_oe : iof0Ctrl_17_oe;
  assign T_8187_ie = T_8186 ? iof1Ctrl_17_ie : iof0Ctrl_17_ie;
  assign T_8191 = iofEnReg_io_q[17];
  assign T_8192_oval = T_8191 ? iofPlusSwPinCtrl_17_oval : swPinCtrl_17_oval;
  assign T_8192_oe = T_8191 ? iofPlusSwPinCtrl_17_oe : swPinCtrl_17_oe;
  assign T_8192_ie = T_8191 ? iofPlusSwPinCtrl_17_ie : swPinCtrl_17_ie;
  assign T_8192_pue = T_8191 ? iofPlusSwPinCtrl_17_pue : swPinCtrl_17_pue;
  assign T_8192_ds = T_8191 ? iofPlusSwPinCtrl_17_ds : swPinCtrl_17_ds;
  assign T_8198 = xorReg[17];
  assign T_8199 = T_8192_oval ^ T_8198;
  assign T_8200 = riseIpReg[17];
  assign T_8201 = riseIeReg[17];
  assign T_8202 = T_8200 & T_8201;
  assign T_8203 = fallIpReg[17];
  assign T_8204 = fallIeReg[17];
  assign T_8205 = T_8203 & T_8204;
  assign T_8206 = T_8202 | T_8205;
  assign T_8207 = highIpReg[17];
  assign T_8208 = highIeReg[17];
  assign T_8209 = T_8207 & T_8208;
  assign T_8210 = T_8206 | T_8209;
  assign T_8211 = lowIpReg[17];
  assign T_8212 = lowIeReg[17];
  assign T_8213 = T_8211 & T_8212;
  assign T_8214 = T_8210 | T_8213;
  assign T_8215 = inSyncReg[17];
  assign T_8217 = pueReg_io_q[18];
  assign T_8218 = portReg[18];
  assign T_8219 = oeReg_io_q[18];
  assign T_8220 = dsReg[18];
  assign T_8221 = ieReg_io_q[18];
  assign GEN_309 = io_port_iof_0_18_o_valid ? io_port_iof_0_18_o_oval : swPinCtrl_18_oval;
  assign GEN_310 = io_port_iof_0_18_o_valid ? io_port_iof_0_18_o_oe : swPinCtrl_18_oe;
  assign GEN_311 = io_port_iof_0_18_o_valid ? io_port_iof_0_18_o_ie : swPinCtrl_18_ie;
  assign GEN_312 = io_port_iof_1_18_o_valid ? io_port_iof_1_18_o_oval : swPinCtrl_18_oval;
  assign GEN_313 = io_port_iof_1_18_o_valid ? io_port_iof_1_18_o_oe : swPinCtrl_18_oe;
  assign GEN_314 = io_port_iof_1_18_o_valid ? io_port_iof_1_18_o_ie : swPinCtrl_18_ie;
  assign T_8222 = iofSelReg[18];
  assign T_8223_oval = T_8222 ? iof1Ctrl_18_oval : iof0Ctrl_18_oval;
  assign T_8223_oe = T_8222 ? iof1Ctrl_18_oe : iof0Ctrl_18_oe;
  assign T_8223_ie = T_8222 ? iof1Ctrl_18_ie : iof0Ctrl_18_ie;
  assign T_8227 = iofEnReg_io_q[18];
  assign T_8228_oval = T_8227 ? iofPlusSwPinCtrl_18_oval : swPinCtrl_18_oval;
  assign T_8228_oe = T_8227 ? iofPlusSwPinCtrl_18_oe : swPinCtrl_18_oe;
  assign T_8228_ie = T_8227 ? iofPlusSwPinCtrl_18_ie : swPinCtrl_18_ie;
  assign T_8228_pue = T_8227 ? iofPlusSwPinCtrl_18_pue : swPinCtrl_18_pue;
  assign T_8228_ds = T_8227 ? iofPlusSwPinCtrl_18_ds : swPinCtrl_18_ds;
  assign T_8234 = xorReg[18];
  assign T_8235 = T_8228_oval ^ T_8234;
  assign T_8236 = riseIpReg[18];
  assign T_8237 = riseIeReg[18];
  assign T_8238 = T_8236 & T_8237;
  assign T_8239 = fallIpReg[18];
  assign T_8240 = fallIeReg[18];
  assign T_8241 = T_8239 & T_8240;
  assign T_8242 = T_8238 | T_8241;
  assign T_8243 = highIpReg[18];
  assign T_8244 = highIeReg[18];
  assign T_8245 = T_8243 & T_8244;
  assign T_8246 = T_8242 | T_8245;
  assign T_8247 = lowIpReg[18];
  assign T_8248 = lowIeReg[18];
  assign T_8249 = T_8247 & T_8248;
  assign T_8250 = T_8246 | T_8249;
  assign T_8251 = inSyncReg[18];
  assign T_8253 = pueReg_io_q[19];
  assign T_8254 = portReg[19];
  assign T_8255 = oeReg_io_q[19];
  assign T_8256 = dsReg[19];
  assign T_8257 = ieReg_io_q[19];
  assign GEN_315 = io_port_iof_0_19_o_valid ? io_port_iof_0_19_o_oval : swPinCtrl_19_oval;
  assign GEN_316 = io_port_iof_0_19_o_valid ? io_port_iof_0_19_o_oe : swPinCtrl_19_oe;
  assign GEN_317 = io_port_iof_0_19_o_valid ? io_port_iof_0_19_o_ie : swPinCtrl_19_ie;
  assign GEN_318 = io_port_iof_1_19_o_valid ? io_port_iof_1_19_o_oval : swPinCtrl_19_oval;
  assign GEN_319 = io_port_iof_1_19_o_valid ? io_port_iof_1_19_o_oe : swPinCtrl_19_oe;
  assign GEN_320 = io_port_iof_1_19_o_valid ? io_port_iof_1_19_o_ie : swPinCtrl_19_ie;
  assign T_8258 = iofSelReg[19];
  assign T_8259_oval = T_8258 ? iof1Ctrl_19_oval : iof0Ctrl_19_oval;
  assign T_8259_oe = T_8258 ? iof1Ctrl_19_oe : iof0Ctrl_19_oe;
  assign T_8259_ie = T_8258 ? iof1Ctrl_19_ie : iof0Ctrl_19_ie;
  assign T_8263 = iofEnReg_io_q[19];
  assign T_8264_oval = T_8263 ? iofPlusSwPinCtrl_19_oval : swPinCtrl_19_oval;
  assign T_8264_oe = T_8263 ? iofPlusSwPinCtrl_19_oe : swPinCtrl_19_oe;
  assign T_8264_ie = T_8263 ? iofPlusSwPinCtrl_19_ie : swPinCtrl_19_ie;
  assign T_8264_pue = T_8263 ? iofPlusSwPinCtrl_19_pue : swPinCtrl_19_pue;
  assign T_8264_ds = T_8263 ? iofPlusSwPinCtrl_19_ds : swPinCtrl_19_ds;
  assign T_8270 = xorReg[19];
  assign T_8271 = T_8264_oval ^ T_8270;
  assign T_8272 = riseIpReg[19];
  assign T_8273 = riseIeReg[19];
  assign T_8274 = T_8272 & T_8273;
  assign T_8275 = fallIpReg[19];
  assign T_8276 = fallIeReg[19];
  assign T_8277 = T_8275 & T_8276;
  assign T_8278 = T_8274 | T_8277;
  assign T_8279 = highIpReg[19];
  assign T_8280 = highIeReg[19];
  assign T_8281 = T_8279 & T_8280;
  assign T_8282 = T_8278 | T_8281;
  assign T_8283 = lowIpReg[19];
  assign T_8284 = lowIeReg[19];
  assign T_8285 = T_8283 & T_8284;
  assign T_8286 = T_8282 | T_8285;
  assign T_8287 = inSyncReg[19];
  assign T_8289 = pueReg_io_q[20];
  assign T_8290 = portReg[20];
  assign T_8291 = oeReg_io_q[20];
  assign T_8292 = dsReg[20];
  assign T_8293 = ieReg_io_q[20];
  assign GEN_321 = io_port_iof_0_20_o_valid ? io_port_iof_0_20_o_oval : swPinCtrl_20_oval;
  assign GEN_322 = io_port_iof_0_20_o_valid ? io_port_iof_0_20_o_oe : swPinCtrl_20_oe;
  assign GEN_323 = io_port_iof_0_20_o_valid ? io_port_iof_0_20_o_ie : swPinCtrl_20_ie;
  assign GEN_324 = io_port_iof_1_20_o_valid ? io_port_iof_1_20_o_oval : swPinCtrl_20_oval;
  assign GEN_325 = io_port_iof_1_20_o_valid ? io_port_iof_1_20_o_oe : swPinCtrl_20_oe;
  assign GEN_326 = io_port_iof_1_20_o_valid ? io_port_iof_1_20_o_ie : swPinCtrl_20_ie;
  assign T_8294 = iofSelReg[20];
  assign T_8295_oval = T_8294 ? iof1Ctrl_20_oval : iof0Ctrl_20_oval;
  assign T_8295_oe = T_8294 ? iof1Ctrl_20_oe : iof0Ctrl_20_oe;
  assign T_8295_ie = T_8294 ? iof1Ctrl_20_ie : iof0Ctrl_20_ie;
  assign T_8299 = iofEnReg_io_q[20];
  assign T_8300_oval = T_8299 ? iofPlusSwPinCtrl_20_oval : swPinCtrl_20_oval;
  assign T_8300_oe = T_8299 ? iofPlusSwPinCtrl_20_oe : swPinCtrl_20_oe;
  assign T_8300_ie = T_8299 ? iofPlusSwPinCtrl_20_ie : swPinCtrl_20_ie;
  assign T_8300_pue = T_8299 ? iofPlusSwPinCtrl_20_pue : swPinCtrl_20_pue;
  assign T_8300_ds = T_8299 ? iofPlusSwPinCtrl_20_ds : swPinCtrl_20_ds;
  assign T_8306 = xorReg[20];
  assign T_8307 = T_8300_oval ^ T_8306;
  assign T_8308 = riseIpReg[20];
  assign T_8309 = riseIeReg[20];
  assign T_8310 = T_8308 & T_8309;
  assign T_8311 = fallIpReg[20];
  assign T_8312 = fallIeReg[20];
  assign T_8313 = T_8311 & T_8312;
  assign T_8314 = T_8310 | T_8313;
  assign T_8315 = highIpReg[20];
  assign T_8316 = highIeReg[20];
  assign T_8317 = T_8315 & T_8316;
  assign T_8318 = T_8314 | T_8317;
  assign T_8319 = lowIpReg[20];
  assign T_8320 = lowIeReg[20];
  assign T_8321 = T_8319 & T_8320;
  assign T_8322 = T_8318 | T_8321;
  assign T_8323 = inSyncReg[20];
  assign T_8325 = pueReg_io_q[21];
  assign T_8326 = portReg[21];
  assign T_8327 = oeReg_io_q[21];
  assign T_8328 = dsReg[21];
  assign T_8329 = ieReg_io_q[21];
  assign GEN_327 = io_port_iof_0_21_o_valid ? io_port_iof_0_21_o_oval : swPinCtrl_21_oval;
  assign GEN_328 = io_port_iof_0_21_o_valid ? io_port_iof_0_21_o_oe : swPinCtrl_21_oe;
  assign GEN_329 = io_port_iof_0_21_o_valid ? io_port_iof_0_21_o_ie : swPinCtrl_21_ie;
  assign GEN_330 = io_port_iof_1_21_o_valid ? io_port_iof_1_21_o_oval : swPinCtrl_21_oval;
  assign GEN_331 = io_port_iof_1_21_o_valid ? io_port_iof_1_21_o_oe : swPinCtrl_21_oe;
  assign GEN_332 = io_port_iof_1_21_o_valid ? io_port_iof_1_21_o_ie : swPinCtrl_21_ie;
  assign T_8330 = iofSelReg[21];
  assign T_8331_oval = T_8330 ? iof1Ctrl_21_oval : iof0Ctrl_21_oval;
  assign T_8331_oe = T_8330 ? iof1Ctrl_21_oe : iof0Ctrl_21_oe;
  assign T_8331_ie = T_8330 ? iof1Ctrl_21_ie : iof0Ctrl_21_ie;
  assign T_8335 = iofEnReg_io_q[21];
  assign T_8336_oval = T_8335 ? iofPlusSwPinCtrl_21_oval : swPinCtrl_21_oval;
  assign T_8336_oe = T_8335 ? iofPlusSwPinCtrl_21_oe : swPinCtrl_21_oe;
  assign T_8336_ie = T_8335 ? iofPlusSwPinCtrl_21_ie : swPinCtrl_21_ie;
  assign T_8336_pue = T_8335 ? iofPlusSwPinCtrl_21_pue : swPinCtrl_21_pue;
  assign T_8336_ds = T_8335 ? iofPlusSwPinCtrl_21_ds : swPinCtrl_21_ds;
  assign T_8342 = xorReg[21];
  assign T_8343 = T_8336_oval ^ T_8342;
  assign T_8344 = riseIpReg[21];
  assign T_8345 = riseIeReg[21];
  assign T_8346 = T_8344 & T_8345;
  assign T_8347 = fallIpReg[21];
  assign T_8348 = fallIeReg[21];
  assign T_8349 = T_8347 & T_8348;
  assign T_8350 = T_8346 | T_8349;
  assign T_8351 = highIpReg[21];
  assign T_8352 = highIeReg[21];
  assign T_8353 = T_8351 & T_8352;
  assign T_8354 = T_8350 | T_8353;
  assign T_8355 = lowIpReg[21];
  assign T_8356 = lowIeReg[21];
  assign T_8357 = T_8355 & T_8356;
  assign T_8358 = T_8354 | T_8357;
  assign T_8359 = inSyncReg[21];
  assign T_8361 = pueReg_io_q[22];
  assign T_8362 = portReg[22];
  assign T_8363 = oeReg_io_q[22];
  assign T_8364 = dsReg[22];
  assign T_8365 = ieReg_io_q[22];
  assign GEN_333 = io_port_iof_0_22_o_valid ? io_port_iof_0_22_o_oval : swPinCtrl_22_oval;
  assign GEN_334 = io_port_iof_0_22_o_valid ? io_port_iof_0_22_o_oe : swPinCtrl_22_oe;
  assign GEN_335 = io_port_iof_0_22_o_valid ? io_port_iof_0_22_o_ie : swPinCtrl_22_ie;
  assign GEN_336 = io_port_iof_1_22_o_valid ? io_port_iof_1_22_o_oval : swPinCtrl_22_oval;
  assign GEN_337 = io_port_iof_1_22_o_valid ? io_port_iof_1_22_o_oe : swPinCtrl_22_oe;
  assign GEN_338 = io_port_iof_1_22_o_valid ? io_port_iof_1_22_o_ie : swPinCtrl_22_ie;
  assign T_8366 = iofSelReg[22];
  assign T_8367_oval = T_8366 ? iof1Ctrl_22_oval : iof0Ctrl_22_oval;
  assign T_8367_oe = T_8366 ? iof1Ctrl_22_oe : iof0Ctrl_22_oe;
  assign T_8367_ie = T_8366 ? iof1Ctrl_22_ie : iof0Ctrl_22_ie;
  assign T_8371 = iofEnReg_io_q[22];
  assign T_8372_oval = T_8371 ? iofPlusSwPinCtrl_22_oval : swPinCtrl_22_oval;
  assign T_8372_oe = T_8371 ? iofPlusSwPinCtrl_22_oe : swPinCtrl_22_oe;
  assign T_8372_ie = T_8371 ? iofPlusSwPinCtrl_22_ie : swPinCtrl_22_ie;
  assign T_8372_pue = T_8371 ? iofPlusSwPinCtrl_22_pue : swPinCtrl_22_pue;
  assign T_8372_ds = T_8371 ? iofPlusSwPinCtrl_22_ds : swPinCtrl_22_ds;
  assign T_8378 = xorReg[22];
  assign T_8379 = T_8372_oval ^ T_8378;
  assign T_8380 = riseIpReg[22];
  assign T_8381 = riseIeReg[22];
  assign T_8382 = T_8380 & T_8381;
  assign T_8383 = fallIpReg[22];
  assign T_8384 = fallIeReg[22];
  assign T_8385 = T_8383 & T_8384;
  assign T_8386 = T_8382 | T_8385;
  assign T_8387 = highIpReg[22];
  assign T_8388 = highIeReg[22];
  assign T_8389 = T_8387 & T_8388;
  assign T_8390 = T_8386 | T_8389;
  assign T_8391 = lowIpReg[22];
  assign T_8392 = lowIeReg[22];
  assign T_8393 = T_8391 & T_8392;
  assign T_8394 = T_8390 | T_8393;
  assign T_8395 = inSyncReg[22];
  assign T_8397 = pueReg_io_q[23];
  assign T_8398 = portReg[23];
  assign T_8399 = oeReg_io_q[23];
  assign T_8400 = dsReg[23];
  assign T_8401 = ieReg_io_q[23];
  assign GEN_339 = io_port_iof_0_23_o_valid ? io_port_iof_0_23_o_oval : swPinCtrl_23_oval;
  assign GEN_340 = io_port_iof_0_23_o_valid ? io_port_iof_0_23_o_oe : swPinCtrl_23_oe;
  assign GEN_341 = io_port_iof_0_23_o_valid ? io_port_iof_0_23_o_ie : swPinCtrl_23_ie;
  assign GEN_342 = io_port_iof_1_23_o_valid ? io_port_iof_1_23_o_oval : swPinCtrl_23_oval;
  assign GEN_343 = io_port_iof_1_23_o_valid ? io_port_iof_1_23_o_oe : swPinCtrl_23_oe;
  assign GEN_344 = io_port_iof_1_23_o_valid ? io_port_iof_1_23_o_ie : swPinCtrl_23_ie;
  assign T_8402 = iofSelReg[23];
  assign T_8403_oval = T_8402 ? iof1Ctrl_23_oval : iof0Ctrl_23_oval;
  assign T_8403_oe = T_8402 ? iof1Ctrl_23_oe : iof0Ctrl_23_oe;
  assign T_8403_ie = T_8402 ? iof1Ctrl_23_ie : iof0Ctrl_23_ie;
  assign T_8407 = iofEnReg_io_q[23];
  assign T_8408_oval = T_8407 ? iofPlusSwPinCtrl_23_oval : swPinCtrl_23_oval;
  assign T_8408_oe = T_8407 ? iofPlusSwPinCtrl_23_oe : swPinCtrl_23_oe;
  assign T_8408_ie = T_8407 ? iofPlusSwPinCtrl_23_ie : swPinCtrl_23_ie;
  assign T_8408_pue = T_8407 ? iofPlusSwPinCtrl_23_pue : swPinCtrl_23_pue;
  assign T_8408_ds = T_8407 ? iofPlusSwPinCtrl_23_ds : swPinCtrl_23_ds;
  assign T_8414 = xorReg[23];
  assign T_8415 = T_8408_oval ^ T_8414;
  assign T_8416 = riseIpReg[23];
  assign T_8417 = riseIeReg[23];
  assign T_8418 = T_8416 & T_8417;
  assign T_8419 = fallIpReg[23];
  assign T_8420 = fallIeReg[23];
  assign T_8421 = T_8419 & T_8420;
  assign T_8422 = T_8418 | T_8421;
  assign T_8423 = highIpReg[23];
  assign T_8424 = highIeReg[23];
  assign T_8425 = T_8423 & T_8424;
  assign T_8426 = T_8422 | T_8425;
  assign T_8427 = lowIpReg[23];
  assign T_8428 = lowIeReg[23];
  assign T_8429 = T_8427 & T_8428;
  assign T_8430 = T_8426 | T_8429;
  assign T_8431 = inSyncReg[23];
  assign T_8433 = pueReg_io_q[24];
  assign T_8434 = portReg[24];
  assign T_8435 = oeReg_io_q[24];
  assign T_8436 = dsReg[24];
  assign T_8437 = ieReg_io_q[24];
  assign GEN_345 = io_port_iof_0_24_o_valid ? io_port_iof_0_24_o_oval : swPinCtrl_24_oval;
  assign GEN_346 = io_port_iof_0_24_o_valid ? io_port_iof_0_24_o_oe : swPinCtrl_24_oe;
  assign GEN_347 = io_port_iof_0_24_o_valid ? io_port_iof_0_24_o_ie : swPinCtrl_24_ie;
  assign GEN_348 = io_port_iof_1_24_o_valid ? io_port_iof_1_24_o_oval : swPinCtrl_24_oval;
  assign GEN_349 = io_port_iof_1_24_o_valid ? io_port_iof_1_24_o_oe : swPinCtrl_24_oe;
  assign GEN_350 = io_port_iof_1_24_o_valid ? io_port_iof_1_24_o_ie : swPinCtrl_24_ie;
  assign T_8438 = iofSelReg[24];
  assign T_8439_oval = T_8438 ? iof1Ctrl_24_oval : iof0Ctrl_24_oval;
  assign T_8439_oe = T_8438 ? iof1Ctrl_24_oe : iof0Ctrl_24_oe;
  assign T_8439_ie = T_8438 ? iof1Ctrl_24_ie : iof0Ctrl_24_ie;
  assign T_8443 = iofEnReg_io_q[24];
  assign T_8444_oval = T_8443 ? iofPlusSwPinCtrl_24_oval : swPinCtrl_24_oval;
  assign T_8444_oe = T_8443 ? iofPlusSwPinCtrl_24_oe : swPinCtrl_24_oe;
  assign T_8444_ie = T_8443 ? iofPlusSwPinCtrl_24_ie : swPinCtrl_24_ie;
  assign T_8444_pue = T_8443 ? iofPlusSwPinCtrl_24_pue : swPinCtrl_24_pue;
  assign T_8444_ds = T_8443 ? iofPlusSwPinCtrl_24_ds : swPinCtrl_24_ds;
  assign T_8450 = xorReg[24];
  assign T_8451 = T_8444_oval ^ T_8450;
  assign T_8452 = riseIpReg[24];
  assign T_8453 = riseIeReg[24];
  assign T_8454 = T_8452 & T_8453;
  assign T_8455 = fallIpReg[24];
  assign T_8456 = fallIeReg[24];
  assign T_8457 = T_8455 & T_8456;
  assign T_8458 = T_8454 | T_8457;
  assign T_8459 = highIpReg[24];
  assign T_8460 = highIeReg[24];
  assign T_8461 = T_8459 & T_8460;
  assign T_8462 = T_8458 | T_8461;
  assign T_8463 = lowIpReg[24];
  assign T_8464 = lowIeReg[24];
  assign T_8465 = T_8463 & T_8464;
  assign T_8466 = T_8462 | T_8465;
  assign T_8467 = inSyncReg[24];
  assign T_8469 = pueReg_io_q[25];
  assign T_8470 = portReg[25];
  assign T_8471 = oeReg_io_q[25];
  assign T_8472 = dsReg[25];
  assign T_8473 = ieReg_io_q[25];
  assign GEN_351 = io_port_iof_0_25_o_valid ? io_port_iof_0_25_o_oval : swPinCtrl_25_oval;
  assign GEN_352 = io_port_iof_0_25_o_valid ? io_port_iof_0_25_o_oe : swPinCtrl_25_oe;
  assign GEN_353 = io_port_iof_0_25_o_valid ? io_port_iof_0_25_o_ie : swPinCtrl_25_ie;
  assign GEN_354 = io_port_iof_1_25_o_valid ? io_port_iof_1_25_o_oval : swPinCtrl_25_oval;
  assign GEN_355 = io_port_iof_1_25_o_valid ? io_port_iof_1_25_o_oe : swPinCtrl_25_oe;
  assign GEN_356 = io_port_iof_1_25_o_valid ? io_port_iof_1_25_o_ie : swPinCtrl_25_ie;
  assign T_8474 = iofSelReg[25];
  assign T_8475_oval = T_8474 ? iof1Ctrl_25_oval : iof0Ctrl_25_oval;
  assign T_8475_oe = T_8474 ? iof1Ctrl_25_oe : iof0Ctrl_25_oe;
  assign T_8475_ie = T_8474 ? iof1Ctrl_25_ie : iof0Ctrl_25_ie;
  assign T_8479 = iofEnReg_io_q[25];
  assign T_8480_oval = T_8479 ? iofPlusSwPinCtrl_25_oval : swPinCtrl_25_oval;
  assign T_8480_oe = T_8479 ? iofPlusSwPinCtrl_25_oe : swPinCtrl_25_oe;
  assign T_8480_ie = T_8479 ? iofPlusSwPinCtrl_25_ie : swPinCtrl_25_ie;
  assign T_8480_pue = T_8479 ? iofPlusSwPinCtrl_25_pue : swPinCtrl_25_pue;
  assign T_8480_ds = T_8479 ? iofPlusSwPinCtrl_25_ds : swPinCtrl_25_ds;
  assign T_8486 = xorReg[25];
  assign T_8487 = T_8480_oval ^ T_8486;
  assign T_8488 = riseIpReg[25];
  assign T_8489 = riseIeReg[25];
  assign T_8490 = T_8488 & T_8489;
  assign T_8491 = fallIpReg[25];
  assign T_8492 = fallIeReg[25];
  assign T_8493 = T_8491 & T_8492;
  assign T_8494 = T_8490 | T_8493;
  assign T_8495 = highIpReg[25];
  assign T_8496 = highIeReg[25];
  assign T_8497 = T_8495 & T_8496;
  assign T_8498 = T_8494 | T_8497;
  assign T_8499 = lowIpReg[25];
  assign T_8500 = lowIeReg[25];
  assign T_8501 = T_8499 & T_8500;
  assign T_8502 = T_8498 | T_8501;
  assign T_8503 = inSyncReg[25];
  assign T_8505 = pueReg_io_q[26];
  assign T_8506 = portReg[26];
  assign T_8507 = oeReg_io_q[26];
  assign T_8508 = dsReg[26];
  assign T_8509 = ieReg_io_q[26];
  assign GEN_357 = io_port_iof_0_26_o_valid ? io_port_iof_0_26_o_oval : swPinCtrl_26_oval;
  assign GEN_358 = io_port_iof_0_26_o_valid ? io_port_iof_0_26_o_oe : swPinCtrl_26_oe;
  assign GEN_359 = io_port_iof_0_26_o_valid ? io_port_iof_0_26_o_ie : swPinCtrl_26_ie;
  assign GEN_360 = io_port_iof_1_26_o_valid ? io_port_iof_1_26_o_oval : swPinCtrl_26_oval;
  assign GEN_361 = io_port_iof_1_26_o_valid ? io_port_iof_1_26_o_oe : swPinCtrl_26_oe;
  assign GEN_362 = io_port_iof_1_26_o_valid ? io_port_iof_1_26_o_ie : swPinCtrl_26_ie;
  assign T_8510 = iofSelReg[26];
  assign T_8511_oval = T_8510 ? iof1Ctrl_26_oval : iof0Ctrl_26_oval;
  assign T_8511_oe = T_8510 ? iof1Ctrl_26_oe : iof0Ctrl_26_oe;
  assign T_8511_ie = T_8510 ? iof1Ctrl_26_ie : iof0Ctrl_26_ie;
  assign T_8515 = iofEnReg_io_q[26];
  assign T_8516_oval = T_8515 ? iofPlusSwPinCtrl_26_oval : swPinCtrl_26_oval;
  assign T_8516_oe = T_8515 ? iofPlusSwPinCtrl_26_oe : swPinCtrl_26_oe;
  assign T_8516_ie = T_8515 ? iofPlusSwPinCtrl_26_ie : swPinCtrl_26_ie;
  assign T_8516_pue = T_8515 ? iofPlusSwPinCtrl_26_pue : swPinCtrl_26_pue;
  assign T_8516_ds = T_8515 ? iofPlusSwPinCtrl_26_ds : swPinCtrl_26_ds;
  assign T_8522 = xorReg[26];
  assign T_8523 = T_8516_oval ^ T_8522;
  assign T_8524 = riseIpReg[26];
  assign T_8525 = riseIeReg[26];
  assign T_8526 = T_8524 & T_8525;
  assign T_8527 = fallIpReg[26];
  assign T_8528 = fallIeReg[26];
  assign T_8529 = T_8527 & T_8528;
  assign T_8530 = T_8526 | T_8529;
  assign T_8531 = highIpReg[26];
  assign T_8532 = highIeReg[26];
  assign T_8533 = T_8531 & T_8532;
  assign T_8534 = T_8530 | T_8533;
  assign T_8535 = lowIpReg[26];
  assign T_8536 = lowIeReg[26];
  assign T_8537 = T_8535 & T_8536;
  assign T_8538 = T_8534 | T_8537;
  assign T_8539 = inSyncReg[26];
  assign T_8541 = pueReg_io_q[27];
  assign T_8542 = portReg[27];
  assign T_8543 = oeReg_io_q[27];
  assign T_8544 = dsReg[27];
  assign T_8545 = ieReg_io_q[27];
  assign GEN_363 = io_port_iof_0_27_o_valid ? io_port_iof_0_27_o_oval : swPinCtrl_27_oval;
  assign GEN_364 = io_port_iof_0_27_o_valid ? io_port_iof_0_27_o_oe : swPinCtrl_27_oe;
  assign GEN_365 = io_port_iof_0_27_o_valid ? io_port_iof_0_27_o_ie : swPinCtrl_27_ie;
  assign GEN_366 = io_port_iof_1_27_o_valid ? io_port_iof_1_27_o_oval : swPinCtrl_27_oval;
  assign GEN_367 = io_port_iof_1_27_o_valid ? io_port_iof_1_27_o_oe : swPinCtrl_27_oe;
  assign GEN_368 = io_port_iof_1_27_o_valid ? io_port_iof_1_27_o_ie : swPinCtrl_27_ie;
  assign T_8546 = iofSelReg[27];
  assign T_8547_oval = T_8546 ? iof1Ctrl_27_oval : iof0Ctrl_27_oval;
  assign T_8547_oe = T_8546 ? iof1Ctrl_27_oe : iof0Ctrl_27_oe;
  assign T_8547_ie = T_8546 ? iof1Ctrl_27_ie : iof0Ctrl_27_ie;
  assign T_8551 = iofEnReg_io_q[27];
  assign T_8552_oval = T_8551 ? iofPlusSwPinCtrl_27_oval : swPinCtrl_27_oval;
  assign T_8552_oe = T_8551 ? iofPlusSwPinCtrl_27_oe : swPinCtrl_27_oe;
  assign T_8552_ie = T_8551 ? iofPlusSwPinCtrl_27_ie : swPinCtrl_27_ie;
  assign T_8552_pue = T_8551 ? iofPlusSwPinCtrl_27_pue : swPinCtrl_27_pue;
  assign T_8552_ds = T_8551 ? iofPlusSwPinCtrl_27_ds : swPinCtrl_27_ds;
  assign T_8558 = xorReg[27];
  assign T_8559 = T_8552_oval ^ T_8558;
  assign T_8560 = riseIpReg[27];
  assign T_8561 = riseIeReg[27];
  assign T_8562 = T_8560 & T_8561;
  assign T_8563 = fallIpReg[27];
  assign T_8564 = fallIeReg[27];
  assign T_8565 = T_8563 & T_8564;
  assign T_8566 = T_8562 | T_8565;
  assign T_8567 = highIpReg[27];
  assign T_8568 = highIeReg[27];
  assign T_8569 = T_8567 & T_8568;
  assign T_8570 = T_8566 | T_8569;
  assign T_8571 = lowIpReg[27];
  assign T_8572 = lowIeReg[27];
  assign T_8573 = T_8571 & T_8572;
  assign T_8574 = T_8570 | T_8573;
  assign T_8575 = inSyncReg[27];
  assign T_8577 = pueReg_io_q[28];
  assign T_8578 = portReg[28];
  assign T_8579 = oeReg_io_q[28];
  assign T_8580 = dsReg[28];
  assign T_8581 = ieReg_io_q[28];
  assign GEN_369 = io_port_iof_0_28_o_valid ? io_port_iof_0_28_o_oval : swPinCtrl_28_oval;
  assign GEN_370 = io_port_iof_0_28_o_valid ? io_port_iof_0_28_o_oe : swPinCtrl_28_oe;
  assign GEN_371 = io_port_iof_0_28_o_valid ? io_port_iof_0_28_o_ie : swPinCtrl_28_ie;
  assign GEN_372 = io_port_iof_1_28_o_valid ? io_port_iof_1_28_o_oval : swPinCtrl_28_oval;
  assign GEN_373 = io_port_iof_1_28_o_valid ? io_port_iof_1_28_o_oe : swPinCtrl_28_oe;
  assign GEN_374 = io_port_iof_1_28_o_valid ? io_port_iof_1_28_o_ie : swPinCtrl_28_ie;
  assign T_8582 = iofSelReg[28];
  assign T_8583_oval = T_8582 ? iof1Ctrl_28_oval : iof0Ctrl_28_oval;
  assign T_8583_oe = T_8582 ? iof1Ctrl_28_oe : iof0Ctrl_28_oe;
  assign T_8583_ie = T_8582 ? iof1Ctrl_28_ie : iof0Ctrl_28_ie;
  assign T_8587 = iofEnReg_io_q[28];
  assign T_8588_oval = T_8587 ? iofPlusSwPinCtrl_28_oval : swPinCtrl_28_oval;
  assign T_8588_oe = T_8587 ? iofPlusSwPinCtrl_28_oe : swPinCtrl_28_oe;
  assign T_8588_ie = T_8587 ? iofPlusSwPinCtrl_28_ie : swPinCtrl_28_ie;
  assign T_8588_pue = T_8587 ? iofPlusSwPinCtrl_28_pue : swPinCtrl_28_pue;
  assign T_8588_ds = T_8587 ? iofPlusSwPinCtrl_28_ds : swPinCtrl_28_ds;
  assign T_8594 = xorReg[28];
  assign T_8595 = T_8588_oval ^ T_8594;
  assign T_8596 = riseIpReg[28];
  assign T_8597 = riseIeReg[28];
  assign T_8598 = T_8596 & T_8597;
  assign T_8599 = fallIpReg[28];
  assign T_8600 = fallIeReg[28];
  assign T_8601 = T_8599 & T_8600;
  assign T_8602 = T_8598 | T_8601;
  assign T_8603 = highIpReg[28];
  assign T_8604 = highIeReg[28];
  assign T_8605 = T_8603 & T_8604;
  assign T_8606 = T_8602 | T_8605;
  assign T_8607 = lowIpReg[28];
  assign T_8608 = lowIeReg[28];
  assign T_8609 = T_8607 & T_8608;
  assign T_8610 = T_8606 | T_8609;
  assign T_8611 = inSyncReg[28];
  assign T_8613 = pueReg_io_q[29];
  assign T_8614 = portReg[29];
  assign T_8615 = oeReg_io_q[29];
  assign T_8616 = dsReg[29];
  assign T_8617 = ieReg_io_q[29];
  assign GEN_375 = io_port_iof_0_29_o_valid ? io_port_iof_0_29_o_oval : swPinCtrl_29_oval;
  assign GEN_376 = io_port_iof_0_29_o_valid ? io_port_iof_0_29_o_oe : swPinCtrl_29_oe;
  assign GEN_377 = io_port_iof_0_29_o_valid ? io_port_iof_0_29_o_ie : swPinCtrl_29_ie;
  assign GEN_378 = io_port_iof_1_29_o_valid ? io_port_iof_1_29_o_oval : swPinCtrl_29_oval;
  assign GEN_379 = io_port_iof_1_29_o_valid ? io_port_iof_1_29_o_oe : swPinCtrl_29_oe;
  assign GEN_380 = io_port_iof_1_29_o_valid ? io_port_iof_1_29_o_ie : swPinCtrl_29_ie;
  assign T_8618 = iofSelReg[29];
  assign T_8619_oval = T_8618 ? iof1Ctrl_29_oval : iof0Ctrl_29_oval;
  assign T_8619_oe = T_8618 ? iof1Ctrl_29_oe : iof0Ctrl_29_oe;
  assign T_8619_ie = T_8618 ? iof1Ctrl_29_ie : iof0Ctrl_29_ie;
  assign T_8623 = iofEnReg_io_q[29];
  assign T_8624_oval = T_8623 ? iofPlusSwPinCtrl_29_oval : swPinCtrl_29_oval;
  assign T_8624_oe = T_8623 ? iofPlusSwPinCtrl_29_oe : swPinCtrl_29_oe;
  assign T_8624_ie = T_8623 ? iofPlusSwPinCtrl_29_ie : swPinCtrl_29_ie;
  assign T_8624_pue = T_8623 ? iofPlusSwPinCtrl_29_pue : swPinCtrl_29_pue;
  assign T_8624_ds = T_8623 ? iofPlusSwPinCtrl_29_ds : swPinCtrl_29_ds;
  assign T_8630 = xorReg[29];
  assign T_8631 = T_8624_oval ^ T_8630;
  assign T_8632 = riseIpReg[29];
  assign T_8633 = riseIeReg[29];
  assign T_8634 = T_8632 & T_8633;
  assign T_8635 = fallIpReg[29];
  assign T_8636 = fallIeReg[29];
  assign T_8637 = T_8635 & T_8636;
  assign T_8638 = T_8634 | T_8637;
  assign T_8639 = highIpReg[29];
  assign T_8640 = highIeReg[29];
  assign T_8641 = T_8639 & T_8640;
  assign T_8642 = T_8638 | T_8641;
  assign T_8643 = lowIpReg[29];
  assign T_8644 = lowIeReg[29];
  assign T_8645 = T_8643 & T_8644;
  assign T_8646 = T_8642 | T_8645;
  assign T_8647 = inSyncReg[29];
  assign T_8649 = pueReg_io_q[30];
  assign T_8650 = portReg[30];
  assign T_8651 = oeReg_io_q[30];
  assign T_8652 = dsReg[30];
  assign T_8653 = ieReg_io_q[30];
  assign GEN_381 = io_port_iof_0_30_o_valid ? io_port_iof_0_30_o_oval : swPinCtrl_30_oval;
  assign GEN_382 = io_port_iof_0_30_o_valid ? io_port_iof_0_30_o_oe : swPinCtrl_30_oe;
  assign GEN_383 = io_port_iof_0_30_o_valid ? io_port_iof_0_30_o_ie : swPinCtrl_30_ie;
  assign GEN_384 = io_port_iof_1_30_o_valid ? io_port_iof_1_30_o_oval : swPinCtrl_30_oval;
  assign GEN_385 = io_port_iof_1_30_o_valid ? io_port_iof_1_30_o_oe : swPinCtrl_30_oe;
  assign GEN_386 = io_port_iof_1_30_o_valid ? io_port_iof_1_30_o_ie : swPinCtrl_30_ie;
  assign T_8654 = iofSelReg[30];
  assign T_8655_oval = T_8654 ? iof1Ctrl_30_oval : iof0Ctrl_30_oval;
  assign T_8655_oe = T_8654 ? iof1Ctrl_30_oe : iof0Ctrl_30_oe;
  assign T_8655_ie = T_8654 ? iof1Ctrl_30_ie : iof0Ctrl_30_ie;
  assign T_8659 = iofEnReg_io_q[30];
  assign T_8660_oval = T_8659 ? iofPlusSwPinCtrl_30_oval : swPinCtrl_30_oval;
  assign T_8660_oe = T_8659 ? iofPlusSwPinCtrl_30_oe : swPinCtrl_30_oe;
  assign T_8660_ie = T_8659 ? iofPlusSwPinCtrl_30_ie : swPinCtrl_30_ie;
  assign T_8660_pue = T_8659 ? iofPlusSwPinCtrl_30_pue : swPinCtrl_30_pue;
  assign T_8660_ds = T_8659 ? iofPlusSwPinCtrl_30_ds : swPinCtrl_30_ds;
  assign T_8666 = xorReg[30];
  assign T_8667 = T_8660_oval ^ T_8666;
  assign T_8668 = riseIpReg[30];
  assign T_8669 = riseIeReg[30];
  assign T_8670 = T_8668 & T_8669;
  assign T_8671 = fallIpReg[30];
  assign T_8672 = fallIeReg[30];
  assign T_8673 = T_8671 & T_8672;
  assign T_8674 = T_8670 | T_8673;
  assign T_8675 = highIpReg[30];
  assign T_8676 = highIeReg[30];
  assign T_8677 = T_8675 & T_8676;
  assign T_8678 = T_8674 | T_8677;
  assign T_8679 = lowIpReg[30];
  assign T_8680 = lowIeReg[30];
  assign T_8681 = T_8679 & T_8680;
  assign T_8682 = T_8678 | T_8681;
  assign T_8683 = inSyncReg[30];
  assign T_8685 = pueReg_io_q[31];
  assign T_8686 = portReg[31];
  assign T_8687 = oeReg_io_q[31];
  assign T_8688 = dsReg[31];
  assign T_8689 = ieReg_io_q[31];
  assign GEN_387 = io_port_iof_0_31_o_valid ? io_port_iof_0_31_o_oval : swPinCtrl_31_oval;
  assign GEN_388 = io_port_iof_0_31_o_valid ? io_port_iof_0_31_o_oe : swPinCtrl_31_oe;
  assign GEN_389 = io_port_iof_0_31_o_valid ? io_port_iof_0_31_o_ie : swPinCtrl_31_ie;
  assign GEN_390 = io_port_iof_1_31_o_valid ? io_port_iof_1_31_o_oval : swPinCtrl_31_oval;
  assign GEN_391 = io_port_iof_1_31_o_valid ? io_port_iof_1_31_o_oe : swPinCtrl_31_oe;
  assign GEN_392 = io_port_iof_1_31_o_valid ? io_port_iof_1_31_o_ie : swPinCtrl_31_ie;
  assign T_8690 = iofSelReg[31];
  assign T_8691_oval = T_8690 ? iof1Ctrl_31_oval : iof0Ctrl_31_oval;
  assign T_8691_oe = T_8690 ? iof1Ctrl_31_oe : iof0Ctrl_31_oe;
  assign T_8691_ie = T_8690 ? iof1Ctrl_31_ie : iof0Ctrl_31_ie;
  assign T_8695 = iofEnReg_io_q[31];
  assign T_8696_oval = T_8695 ? iofPlusSwPinCtrl_31_oval : swPinCtrl_31_oval;
  assign T_8696_oe = T_8695 ? iofPlusSwPinCtrl_31_oe : swPinCtrl_31_oe;
  assign T_8696_ie = T_8695 ? iofPlusSwPinCtrl_31_ie : swPinCtrl_31_ie;
  assign T_8696_pue = T_8695 ? iofPlusSwPinCtrl_31_pue : swPinCtrl_31_pue;
  assign T_8696_ds = T_8695 ? iofPlusSwPinCtrl_31_ds : swPinCtrl_31_ds;
  assign T_8702 = xorReg[31];
  assign T_8703 = T_8696_oval ^ T_8702;
  assign T_8704 = riseIpReg[31];
  assign T_8705 = riseIeReg[31];
  assign T_8706 = T_8704 & T_8705;
  assign T_8707 = fallIpReg[31];
  assign T_8708 = fallIeReg[31];
  assign T_8709 = T_8707 & T_8708;
  assign T_8710 = T_8706 | T_8709;
  assign T_8711 = highIpReg[31];
  assign T_8712 = highIeReg[31];
  assign T_8713 = T_8711 & T_8712;
  assign T_8714 = T_8710 | T_8713;
  assign T_8715 = lowIpReg[31];
  assign T_8716 = lowIeReg[31];
  assign T_8717 = T_8715 & T_8716;
  assign T_8718 = T_8714 | T_8717;
  assign T_8719 = inSyncReg[31];

  always @(posedge clock or posedge reset)
    if(reset) begin
      T_3256 <= 32'b0;
      T_3257 <= 32'b0;
      inSyncReg <= 32'b0;
    end
    else begin
      T_3256 <= inVal;
      T_3257 <= T_3256;
      inSyncReg <= T_3257;
    end

  always @(posedge clock or posedge reset) 
    if (reset) begin
      portReg <= 32'h0;
    end else begin
      if (T_4329) begin
        portReg <= T_3370_bits_data;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      dsReg <= 32'h0;
    end else begin
      if (T_3911) begin
        dsReg <= T_3370_bits_data;
      end
    end


  always @(posedge clock or posedge reset)
    if (reset) begin
      valueReg <= 32'h0;
    end else begin
      valueReg <= inSyncReg;
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      highIeReg <= 32'h0;
    end else begin
      if (T_3951) begin
        highIeReg <= T_3370_bits_data;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      lowIeReg <= 32'h0;
    end else begin
      if (T_4243) begin
        lowIeReg <= T_3370_bits_data;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      riseIeReg <= 32'h0;
    end else begin
      if (T_4071) begin
        riseIeReg <= T_3370_bits_data;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      fallIeReg <= 32'h0;
    end else begin
      if (T_4455) begin
        fallIeReg <= T_3370_bits_data;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      highIpReg <= 32'h0;
    end else begin
      highIpReg <= T_4417;
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      lowIpReg <= 32'h0;
    end else begin
      lowIpReg <= T_4165;
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      riseIpReg <= 32'h0;
    end else begin
      riseIpReg <= T_4291;
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      fallIpReg <= 32'h0;
    end else begin
      fallIpReg <= T_4119;
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      iofSelReg <= 32'h0;
    end else begin
      if (T_4535) begin
        iofSelReg <= T_3370_bits_data;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      xorReg <= 32'h0;
    end else begin
      if (T_4369) begin
        xorReg <= T_3370_bits_data;
      end
    end

endmodule
