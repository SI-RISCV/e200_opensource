 /*                                                                      
 Copyright 2017 Silicon Integrated Microelectronics, Inc.                
                                                                         
 Licensed under the Apache License, Version 2.0 (the "License");         
 you may not use this file except in compliance with the License.        
 You may obtain a copy of the License at                                 
                                                                         
     http://www.apache.org/licenses/LICENSE-2.0                          
                                                                         
  Unless required by applicable law or agreed to in writing, software    
 distributed under the License is distributed on an "AS IS" BASIS,       
 WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 See the License for the specific language governing permissions and     
 limitations under the License.                                          
 */                                                                      
                                                                         
                                                                         
                                                                         

module sirv_plic(
  input   clock,
  input   reset,
  output  io_tl_in_0_a_ready,
  input   io_tl_in_0_a_valid,
  input  [2:0] io_tl_in_0_a_bits_opcode,
  input  [2:0] io_tl_in_0_a_bits_param,
  input  [2:0] io_tl_in_0_a_bits_size,
  input  [4:0] io_tl_in_0_a_bits_source,
  input  [27:0] io_tl_in_0_a_bits_address,
  input  [3:0] io_tl_in_0_a_bits_mask,
  input  [31:0] io_tl_in_0_a_bits_data,
  input   io_tl_in_0_b_ready,
  output  io_tl_in_0_b_valid,
  output [2:0] io_tl_in_0_b_bits_opcode,
  output [1:0] io_tl_in_0_b_bits_param,
  output [2:0] io_tl_in_0_b_bits_size,
  output [4:0] io_tl_in_0_b_bits_source,
  output [27:0] io_tl_in_0_b_bits_address,
  output [3:0] io_tl_in_0_b_bits_mask,
  output [31:0] io_tl_in_0_b_bits_data,
  output  io_tl_in_0_c_ready,
  input   io_tl_in_0_c_valid,
  input  [2:0] io_tl_in_0_c_bits_opcode,
  input  [2:0] io_tl_in_0_c_bits_param,
  input  [2:0] io_tl_in_0_c_bits_size,
  input  [4:0] io_tl_in_0_c_bits_source,
  input  [27:0] io_tl_in_0_c_bits_address,
  input  [31:0] io_tl_in_0_c_bits_data,
  input   io_tl_in_0_c_bits_error,
  input   io_tl_in_0_d_ready,
  output  io_tl_in_0_d_valid,
  output [2:0] io_tl_in_0_d_bits_opcode,
  output [1:0] io_tl_in_0_d_bits_param,
  output [2:0] io_tl_in_0_d_bits_size,
  output [4:0] io_tl_in_0_d_bits_source,
  output  io_tl_in_0_d_bits_sink,
  output [1:0] io_tl_in_0_d_bits_addr_lo,
  output [31:0] io_tl_in_0_d_bits_data,
  output  io_tl_in_0_d_bits_error,
  output  io_tl_in_0_e_ready,
  input   io_tl_in_0_e_valid,
  input   io_tl_in_0_e_bits_sink,
  input   io_devices_0_0,
  input   io_devices_0_1,
  input   io_devices_0_2,
  input   io_devices_0_3,
  input   io_devices_0_4,
  input   io_devices_0_5,
  input   io_devices_0_6,
  input   io_devices_0_7,
  input   io_devices_0_8,
  input   io_devices_0_9,
  input   io_devices_0_10,
  input   io_devices_0_11,
  input   io_devices_0_12,
  input   io_devices_0_13,
  input   io_devices_0_14,
  input   io_devices_0_15,
  input   io_devices_0_16,
  input   io_devices_0_17,
  input   io_devices_0_18,
  input   io_devices_0_19,
  input   io_devices_0_20,
  input   io_devices_0_21,
  input   io_devices_0_22,
  input   io_devices_0_23,
  input   io_devices_0_24,
  input   io_devices_0_25,
  input   io_devices_0_26,
  input   io_devices_0_27,
  input   io_devices_0_28,
  input   io_devices_0_29,
  input   io_devices_0_30,
  input   io_devices_0_31,
  input   io_devices_0_32,
  input   io_devices_0_33,
  input   io_devices_0_34,
  input   io_devices_0_35,
  input   io_devices_0_36,
  input   io_devices_0_37,
  input   io_devices_0_38,
  input   io_devices_0_39,
  input   io_devices_0_40,
  input   io_devices_0_41,
  input   io_devices_0_42,
  input   io_devices_0_43,
  input   io_devices_0_44,
  input   io_devices_0_45,
  input   io_devices_0_46,
  input   io_devices_0_47,
  input   io_devices_0_48,
  input   io_devices_0_49,
  input   io_devices_0_50,
  output  io_harts_0_0
);
  wire  LevelGateway_51_clock;
  wire  LevelGateway_51_reset;
  wire  LevelGateway_51_io_interrupt;
  wire  LevelGateway_51_io_plic_valid;
  wire  LevelGateway_51_io_plic_ready;
  wire  LevelGateway_51_io_plic_complete;
  wire  LevelGateway_1_1_clock;
  wire  LevelGateway_1_1_reset;
  wire  LevelGateway_1_1_io_interrupt;
  wire  LevelGateway_1_1_io_plic_valid;
  wire  LevelGateway_1_1_io_plic_ready;
  wire  LevelGateway_1_1_io_plic_complete;
  wire  LevelGateway_2_1_clock;
  wire  LevelGateway_2_1_reset;
  wire  LevelGateway_2_1_io_interrupt;
  wire  LevelGateway_2_1_io_plic_valid;
  wire  LevelGateway_2_1_io_plic_ready;
  wire  LevelGateway_2_1_io_plic_complete;
  wire  LevelGateway_3_1_clock;
  wire  LevelGateway_3_1_reset;
  wire  LevelGateway_3_1_io_interrupt;
  wire  LevelGateway_3_1_io_plic_valid;
  wire  LevelGateway_3_1_io_plic_ready;
  wire  LevelGateway_3_1_io_plic_complete;
  wire  LevelGateway_4_1_clock;
  wire  LevelGateway_4_1_reset;
  wire  LevelGateway_4_1_io_interrupt;
  wire  LevelGateway_4_1_io_plic_valid;
  wire  LevelGateway_4_1_io_plic_ready;
  wire  LevelGateway_4_1_io_plic_complete;
  wire  LevelGateway_5_1_clock;
  wire  LevelGateway_5_1_reset;
  wire  LevelGateway_5_1_io_interrupt;
  wire  LevelGateway_5_1_io_plic_valid;
  wire  LevelGateway_5_1_io_plic_ready;
  wire  LevelGateway_5_1_io_plic_complete;
  wire  LevelGateway_6_1_clock;
  wire  LevelGateway_6_1_reset;
  wire  LevelGateway_6_1_io_interrupt;
  wire  LevelGateway_6_1_io_plic_valid;
  wire  LevelGateway_6_1_io_plic_ready;
  wire  LevelGateway_6_1_io_plic_complete;
  wire  LevelGateway_7_1_clock;
  wire  LevelGateway_7_1_reset;
  wire  LevelGateway_7_1_io_interrupt;
  wire  LevelGateway_7_1_io_plic_valid;
  wire  LevelGateway_7_1_io_plic_ready;
  wire  LevelGateway_7_1_io_plic_complete;
  wire  LevelGateway_8_1_clock;
  wire  LevelGateway_8_1_reset;
  wire  LevelGateway_8_1_io_interrupt;
  wire  LevelGateway_8_1_io_plic_valid;
  wire  LevelGateway_8_1_io_plic_ready;
  wire  LevelGateway_8_1_io_plic_complete;
  wire  LevelGateway_9_1_clock;
  wire  LevelGateway_9_1_reset;
  wire  LevelGateway_9_1_io_interrupt;
  wire  LevelGateway_9_1_io_plic_valid;
  wire  LevelGateway_9_1_io_plic_ready;
  wire  LevelGateway_9_1_io_plic_complete;
  wire  LevelGateway_10_1_clock;
  wire  LevelGateway_10_1_reset;
  wire  LevelGateway_10_1_io_interrupt;
  wire  LevelGateway_10_1_io_plic_valid;
  wire  LevelGateway_10_1_io_plic_ready;
  wire  LevelGateway_10_1_io_plic_complete;
  wire  LevelGateway_11_1_clock;
  wire  LevelGateway_11_1_reset;
  wire  LevelGateway_11_1_io_interrupt;
  wire  LevelGateway_11_1_io_plic_valid;
  wire  LevelGateway_11_1_io_plic_ready;
  wire  LevelGateway_11_1_io_plic_complete;
  wire  LevelGateway_12_1_clock;
  wire  LevelGateway_12_1_reset;
  wire  LevelGateway_12_1_io_interrupt;
  wire  LevelGateway_12_1_io_plic_valid;
  wire  LevelGateway_12_1_io_plic_ready;
  wire  LevelGateway_12_1_io_plic_complete;
  wire  LevelGateway_13_1_clock;
  wire  LevelGateway_13_1_reset;
  wire  LevelGateway_13_1_io_interrupt;
  wire  LevelGateway_13_1_io_plic_valid;
  wire  LevelGateway_13_1_io_plic_ready;
  wire  LevelGateway_13_1_io_plic_complete;
  wire  LevelGateway_14_1_clock;
  wire  LevelGateway_14_1_reset;
  wire  LevelGateway_14_1_io_interrupt;
  wire  LevelGateway_14_1_io_plic_valid;
  wire  LevelGateway_14_1_io_plic_ready;
  wire  LevelGateway_14_1_io_plic_complete;
  wire  LevelGateway_15_1_clock;
  wire  LevelGateway_15_1_reset;
  wire  LevelGateway_15_1_io_interrupt;
  wire  LevelGateway_15_1_io_plic_valid;
  wire  LevelGateway_15_1_io_plic_ready;
  wire  LevelGateway_15_1_io_plic_complete;
  wire  LevelGateway_16_1_clock;
  wire  LevelGateway_16_1_reset;
  wire  LevelGateway_16_1_io_interrupt;
  wire  LevelGateway_16_1_io_plic_valid;
  wire  LevelGateway_16_1_io_plic_ready;
  wire  LevelGateway_16_1_io_plic_complete;
  wire  LevelGateway_17_1_clock;
  wire  LevelGateway_17_1_reset;
  wire  LevelGateway_17_1_io_interrupt;
  wire  LevelGateway_17_1_io_plic_valid;
  wire  LevelGateway_17_1_io_plic_ready;
  wire  LevelGateway_17_1_io_plic_complete;
  wire  LevelGateway_18_1_clock;
  wire  LevelGateway_18_1_reset;
  wire  LevelGateway_18_1_io_interrupt;
  wire  LevelGateway_18_1_io_plic_valid;
  wire  LevelGateway_18_1_io_plic_ready;
  wire  LevelGateway_18_1_io_plic_complete;
  wire  LevelGateway_19_1_clock;
  wire  LevelGateway_19_1_reset;
  wire  LevelGateway_19_1_io_interrupt;
  wire  LevelGateway_19_1_io_plic_valid;
  wire  LevelGateway_19_1_io_plic_ready;
  wire  LevelGateway_19_1_io_plic_complete;
  wire  LevelGateway_20_1_clock;
  wire  LevelGateway_20_1_reset;
  wire  LevelGateway_20_1_io_interrupt;
  wire  LevelGateway_20_1_io_plic_valid;
  wire  LevelGateway_20_1_io_plic_ready;
  wire  LevelGateway_20_1_io_plic_complete;
  wire  LevelGateway_21_1_clock;
  wire  LevelGateway_21_1_reset;
  wire  LevelGateway_21_1_io_interrupt;
  wire  LevelGateway_21_1_io_plic_valid;
  wire  LevelGateway_21_1_io_plic_ready;
  wire  LevelGateway_21_1_io_plic_complete;
  wire  LevelGateway_22_1_clock;
  wire  LevelGateway_22_1_reset;
  wire  LevelGateway_22_1_io_interrupt;
  wire  LevelGateway_22_1_io_plic_valid;
  wire  LevelGateway_22_1_io_plic_ready;
  wire  LevelGateway_22_1_io_plic_complete;
  wire  LevelGateway_23_1_clock;
  wire  LevelGateway_23_1_reset;
  wire  LevelGateway_23_1_io_interrupt;
  wire  LevelGateway_23_1_io_plic_valid;
  wire  LevelGateway_23_1_io_plic_ready;
  wire  LevelGateway_23_1_io_plic_complete;
  wire  LevelGateway_24_1_clock;
  wire  LevelGateway_24_1_reset;
  wire  LevelGateway_24_1_io_interrupt;
  wire  LevelGateway_24_1_io_plic_valid;
  wire  LevelGateway_24_1_io_plic_ready;
  wire  LevelGateway_24_1_io_plic_complete;
  wire  LevelGateway_25_1_clock;
  wire  LevelGateway_25_1_reset;
  wire  LevelGateway_25_1_io_interrupt;
  wire  LevelGateway_25_1_io_plic_valid;
  wire  LevelGateway_25_1_io_plic_ready;
  wire  LevelGateway_25_1_io_plic_complete;
  wire  LevelGateway_26_1_clock;
  wire  LevelGateway_26_1_reset;
  wire  LevelGateway_26_1_io_interrupt;
  wire  LevelGateway_26_1_io_plic_valid;
  wire  LevelGateway_26_1_io_plic_ready;
  wire  LevelGateway_26_1_io_plic_complete;
  wire  LevelGateway_27_1_clock;
  wire  LevelGateway_27_1_reset;
  wire  LevelGateway_27_1_io_interrupt;
  wire  LevelGateway_27_1_io_plic_valid;
  wire  LevelGateway_27_1_io_plic_ready;
  wire  LevelGateway_27_1_io_plic_complete;
  wire  LevelGateway_28_1_clock;
  wire  LevelGateway_28_1_reset;
  wire  LevelGateway_28_1_io_interrupt;
  wire  LevelGateway_28_1_io_plic_valid;
  wire  LevelGateway_28_1_io_plic_ready;
  wire  LevelGateway_28_1_io_plic_complete;
  wire  LevelGateway_29_1_clock;
  wire  LevelGateway_29_1_reset;
  wire  LevelGateway_29_1_io_interrupt;
  wire  LevelGateway_29_1_io_plic_valid;
  wire  LevelGateway_29_1_io_plic_ready;
  wire  LevelGateway_29_1_io_plic_complete;
  wire  LevelGateway_30_1_clock;
  wire  LevelGateway_30_1_reset;
  wire  LevelGateway_30_1_io_interrupt;
  wire  LevelGateway_30_1_io_plic_valid;
  wire  LevelGateway_30_1_io_plic_ready;
  wire  LevelGateway_30_1_io_plic_complete;
  wire  LevelGateway_31_1_clock;
  wire  LevelGateway_31_1_reset;
  wire  LevelGateway_31_1_io_interrupt;
  wire  LevelGateway_31_1_io_plic_valid;
  wire  LevelGateway_31_1_io_plic_ready;
  wire  LevelGateway_31_1_io_plic_complete;
  wire  LevelGateway_32_1_clock;
  wire  LevelGateway_32_1_reset;
  wire  LevelGateway_32_1_io_interrupt;
  wire  LevelGateway_32_1_io_plic_valid;
  wire  LevelGateway_32_1_io_plic_ready;
  wire  LevelGateway_32_1_io_plic_complete;
  wire  LevelGateway_33_1_clock;
  wire  LevelGateway_33_1_reset;
  wire  LevelGateway_33_1_io_interrupt;
  wire  LevelGateway_33_1_io_plic_valid;
  wire  LevelGateway_33_1_io_plic_ready;
  wire  LevelGateway_33_1_io_plic_complete;
  wire  LevelGateway_34_1_clock;
  wire  LevelGateway_34_1_reset;
  wire  LevelGateway_34_1_io_interrupt;
  wire  LevelGateway_34_1_io_plic_valid;
  wire  LevelGateway_34_1_io_plic_ready;
  wire  LevelGateway_34_1_io_plic_complete;
  wire  LevelGateway_35_1_clock;
  wire  LevelGateway_35_1_reset;
  wire  LevelGateway_35_1_io_interrupt;
  wire  LevelGateway_35_1_io_plic_valid;
  wire  LevelGateway_35_1_io_plic_ready;
  wire  LevelGateway_35_1_io_plic_complete;
  wire  LevelGateway_36_1_clock;
  wire  LevelGateway_36_1_reset;
  wire  LevelGateway_36_1_io_interrupt;
  wire  LevelGateway_36_1_io_plic_valid;
  wire  LevelGateway_36_1_io_plic_ready;
  wire  LevelGateway_36_1_io_plic_complete;
  wire  LevelGateway_37_1_clock;
  wire  LevelGateway_37_1_reset;
  wire  LevelGateway_37_1_io_interrupt;
  wire  LevelGateway_37_1_io_plic_valid;
  wire  LevelGateway_37_1_io_plic_ready;
  wire  LevelGateway_37_1_io_plic_complete;
  wire  LevelGateway_38_1_clock;
  wire  LevelGateway_38_1_reset;
  wire  LevelGateway_38_1_io_interrupt;
  wire  LevelGateway_38_1_io_plic_valid;
  wire  LevelGateway_38_1_io_plic_ready;
  wire  LevelGateway_38_1_io_plic_complete;
  wire  LevelGateway_39_1_clock;
  wire  LevelGateway_39_1_reset;
  wire  LevelGateway_39_1_io_interrupt;
  wire  LevelGateway_39_1_io_plic_valid;
  wire  LevelGateway_39_1_io_plic_ready;
  wire  LevelGateway_39_1_io_plic_complete;
  wire  LevelGateway_40_1_clock;
  wire  LevelGateway_40_1_reset;
  wire  LevelGateway_40_1_io_interrupt;
  wire  LevelGateway_40_1_io_plic_valid;
  wire  LevelGateway_40_1_io_plic_ready;
  wire  LevelGateway_40_1_io_plic_complete;
  wire  LevelGateway_41_1_clock;
  wire  LevelGateway_41_1_reset;
  wire  LevelGateway_41_1_io_interrupt;
  wire  LevelGateway_41_1_io_plic_valid;
  wire  LevelGateway_41_1_io_plic_ready;
  wire  LevelGateway_41_1_io_plic_complete;
  wire  LevelGateway_42_1_clock;
  wire  LevelGateway_42_1_reset;
  wire  LevelGateway_42_1_io_interrupt;
  wire  LevelGateway_42_1_io_plic_valid;
  wire  LevelGateway_42_1_io_plic_ready;
  wire  LevelGateway_42_1_io_plic_complete;
  wire  LevelGateway_43_1_clock;
  wire  LevelGateway_43_1_reset;
  wire  LevelGateway_43_1_io_interrupt;
  wire  LevelGateway_43_1_io_plic_valid;
  wire  LevelGateway_43_1_io_plic_ready;
  wire  LevelGateway_43_1_io_plic_complete;
  wire  LevelGateway_44_1_clock;
  wire  LevelGateway_44_1_reset;
  wire  LevelGateway_44_1_io_interrupt;
  wire  LevelGateway_44_1_io_plic_valid;
  wire  LevelGateway_44_1_io_plic_ready;
  wire  LevelGateway_44_1_io_plic_complete;
  wire  LevelGateway_45_1_clock;
  wire  LevelGateway_45_1_reset;
  wire  LevelGateway_45_1_io_interrupt;
  wire  LevelGateway_45_1_io_plic_valid;
  wire  LevelGateway_45_1_io_plic_ready;
  wire  LevelGateway_45_1_io_plic_complete;
  wire  LevelGateway_46_1_clock;
  wire  LevelGateway_46_1_reset;
  wire  LevelGateway_46_1_io_interrupt;
  wire  LevelGateway_46_1_io_plic_valid;
  wire  LevelGateway_46_1_io_plic_ready;
  wire  LevelGateway_46_1_io_plic_complete;
  wire  LevelGateway_47_1_clock;
  wire  LevelGateway_47_1_reset;
  wire  LevelGateway_47_1_io_interrupt;
  wire  LevelGateway_47_1_io_plic_valid;
  wire  LevelGateway_47_1_io_plic_ready;
  wire  LevelGateway_47_1_io_plic_complete;
  wire  LevelGateway_48_1_clock;
  wire  LevelGateway_48_1_reset;
  wire  LevelGateway_48_1_io_interrupt;
  wire  LevelGateway_48_1_io_plic_valid;
  wire  LevelGateway_48_1_io_plic_ready;
  wire  LevelGateway_48_1_io_plic_complete;
  wire  LevelGateway_49_1_clock;
  wire  LevelGateway_49_1_reset;
  wire  LevelGateway_49_1_io_interrupt;
  wire  LevelGateway_49_1_io_plic_valid;
  wire  LevelGateway_49_1_io_plic_ready;
  wire  LevelGateway_49_1_io_plic_complete;
  wire  LevelGateway_50_1_clock;
  wire  LevelGateway_50_1_reset;
  wire  LevelGateway_50_1_io_interrupt;
  wire  LevelGateway_50_1_io_plic_valid;
  wire  LevelGateway_50_1_io_plic_ready;
  wire  LevelGateway_50_1_io_plic_complete;
  wire  gateways_0_valid;
  wire  gateways_0_ready;
  wire  gateways_0_complete;
  wire  gateways_1_valid;
  wire  gateways_1_ready;
  wire  gateways_1_complete;
  wire  gateways_2_valid;
  wire  gateways_2_ready;
  wire  gateways_2_complete;
  wire  gateways_3_valid;
  wire  gateways_3_ready;
  wire  gateways_3_complete;
  wire  gateways_4_valid;
  wire  gateways_4_ready;
  wire  gateways_4_complete;
  wire  gateways_5_valid;
  wire  gateways_5_ready;
  wire  gateways_5_complete;
  wire  gateways_6_valid;
  wire  gateways_6_ready;
  wire  gateways_6_complete;
  wire  gateways_7_valid;
  wire  gateways_7_ready;
  wire  gateways_7_complete;
  wire  gateways_8_valid;
  wire  gateways_8_ready;
  wire  gateways_8_complete;
  wire  gateways_9_valid;
  wire  gateways_9_ready;
  wire  gateways_9_complete;
  wire  gateways_10_valid;
  wire  gateways_10_ready;
  wire  gateways_10_complete;
  wire  gateways_11_valid;
  wire  gateways_11_ready;
  wire  gateways_11_complete;
  wire  gateways_12_valid;
  wire  gateways_12_ready;
  wire  gateways_12_complete;
  wire  gateways_13_valid;
  wire  gateways_13_ready;
  wire  gateways_13_complete;
  wire  gateways_14_valid;
  wire  gateways_14_ready;
  wire  gateways_14_complete;
  wire  gateways_15_valid;
  wire  gateways_15_ready;
  wire  gateways_15_complete;
  wire  gateways_16_valid;
  wire  gateways_16_ready;
  wire  gateways_16_complete;
  wire  gateways_17_valid;
  wire  gateways_17_ready;
  wire  gateways_17_complete;
  wire  gateways_18_valid;
  wire  gateways_18_ready;
  wire  gateways_18_complete;
  wire  gateways_19_valid;
  wire  gateways_19_ready;
  wire  gateways_19_complete;
  wire  gateways_20_valid;
  wire  gateways_20_ready;
  wire  gateways_20_complete;
  wire  gateways_21_valid;
  wire  gateways_21_ready;
  wire  gateways_21_complete;
  wire  gateways_22_valid;
  wire  gateways_22_ready;
  wire  gateways_22_complete;
  wire  gateways_23_valid;
  wire  gateways_23_ready;
  wire  gateways_23_complete;
  wire  gateways_24_valid;
  wire  gateways_24_ready;
  wire  gateways_24_complete;
  wire  gateways_25_valid;
  wire  gateways_25_ready;
  wire  gateways_25_complete;
  wire  gateways_26_valid;
  wire  gateways_26_ready;
  wire  gateways_26_complete;
  wire  gateways_27_valid;
  wire  gateways_27_ready;
  wire  gateways_27_complete;
  wire  gateways_28_valid;
  wire  gateways_28_ready;
  wire  gateways_28_complete;
  wire  gateways_29_valid;
  wire  gateways_29_ready;
  wire  gateways_29_complete;
  wire  gateways_30_valid;
  wire  gateways_30_ready;
  wire  gateways_30_complete;
  wire  gateways_31_valid;
  wire  gateways_31_ready;
  wire  gateways_31_complete;
  wire  gateways_32_valid;
  wire  gateways_32_ready;
  wire  gateways_32_complete;
  wire  gateways_33_valid;
  wire  gateways_33_ready;
  wire  gateways_33_complete;
  wire  gateways_34_valid;
  wire  gateways_34_ready;
  wire  gateways_34_complete;
  wire  gateways_35_valid;
  wire  gateways_35_ready;
  wire  gateways_35_complete;
  wire  gateways_36_valid;
  wire  gateways_36_ready;
  wire  gateways_36_complete;
  wire  gateways_37_valid;
  wire  gateways_37_ready;
  wire  gateways_37_complete;
  wire  gateways_38_valid;
  wire  gateways_38_ready;
  wire  gateways_38_complete;
  wire  gateways_39_valid;
  wire  gateways_39_ready;
  wire  gateways_39_complete;
  wire  gateways_40_valid;
  wire  gateways_40_ready;
  wire  gateways_40_complete;
  wire  gateways_41_valid;
  wire  gateways_41_ready;
  wire  gateways_41_complete;
  wire  gateways_42_valid;
  wire  gateways_42_ready;
  wire  gateways_42_complete;
  wire  gateways_43_valid;
  wire  gateways_43_ready;
  wire  gateways_43_complete;
  wire  gateways_44_valid;
  wire  gateways_44_ready;
  wire  gateways_44_complete;
  wire  gateways_45_valid;
  wire  gateways_45_ready;
  wire  gateways_45_complete;
  wire  gateways_46_valid;
  wire  gateways_46_ready;
  wire  gateways_46_complete;
  wire  gateways_47_valid;
  wire  gateways_47_ready;
  wire  gateways_47_complete;
  wire  gateways_48_valid;
  wire  gateways_48_ready;
  wire  gateways_48_complete;
  wire  gateways_49_valid;
  wire  gateways_49_ready;
  wire  gateways_49_complete;
  wire  gateways_50_valid;
  wire  gateways_50_ready;
  wire  gateways_50_complete;
  reg [2:0] priority_0;
  reg [31:0] GEN_3717;
  reg [2:0] priority_1;
  reg [31:0] GEN_3718;
  reg [2:0] priority_2;
  reg [31:0] GEN_3719;
  reg [2:0] priority_3;
  reg [31:0] GEN_3720;
  reg [2:0] priority_4;
  reg [31:0] GEN_3721;
  reg [2:0] priority_5;
  reg [31:0] GEN_3722;
  reg [2:0] priority_6;
  reg [31:0] GEN_3723;
  reg [2:0] priority_7;
  reg [31:0] GEN_3724;
  reg [2:0] priority_8;
  reg [31:0] GEN_3725;
  reg [2:0] priority_9;
  reg [31:0] GEN_3726;
  reg [2:0] priority_10;
  reg [31:0] GEN_3727;
  reg [2:0] priority_11;
  reg [31:0] GEN_3728;
  reg [2:0] priority_12;
  reg [31:0] GEN_3729;
  reg [2:0] priority_13;
  reg [31:0] GEN_3730;
  reg [2:0] priority_14;
  reg [31:0] GEN_3731;
  reg [2:0] priority_15;
  reg [31:0] GEN_3732;
  reg [2:0] priority_16;
  reg [31:0] GEN_3733;
  reg [2:0] priority_17;
  reg [31:0] GEN_3734;
  reg [2:0] priority_18;
  reg [31:0] GEN_3735;
  reg [2:0] priority_19;
  reg [31:0] GEN_3736;
  reg [2:0] priority_20;
  reg [31:0] GEN_3737;
  reg [2:0] priority_21;
  reg [31:0] GEN_3738;
  reg [2:0] priority_22;
  reg [31:0] GEN_3739;
  reg [2:0] priority_23;
  reg [31:0] GEN_3740;
  reg [2:0] priority_24;
  reg [31:0] GEN_3741;
  reg [2:0] priority_25;
  reg [31:0] GEN_3742;
  reg [2:0] priority_26;
  reg [31:0] GEN_3743;
  reg [2:0] priority_27;
  reg [31:0] GEN_3744;
  reg [2:0] priority_28;
  reg [31:0] GEN_3745;
  reg [2:0] priority_29;
  reg [31:0] GEN_3746;
  reg [2:0] priority_30;
  reg [31:0] GEN_3747;
  reg [2:0] priority_31;
  reg [31:0] GEN_3748;
  reg [2:0] priority_32;
  reg [31:0] GEN_3749;
  reg [2:0] priority_33;
  reg [31:0] GEN_3750;
  reg [2:0] priority_34;
  reg [31:0] GEN_3751;
  reg [2:0] priority_35;
  reg [31:0] GEN_3752;
  reg [2:0] priority_36;
  reg [31:0] GEN_3753;
  reg [2:0] priority_37;
  reg [31:0] GEN_3754;
  reg [2:0] priority_38;
  reg [31:0] GEN_3755;
  reg [2:0] priority_39;
  reg [31:0] GEN_3756;
  reg [2:0] priority_40;
  reg [31:0] GEN_3757;
  reg [2:0] priority_41;
  reg [31:0] GEN_3758;
  reg [2:0] priority_42;
  reg [31:0] GEN_3759;
  reg [2:0] priority_43;
  reg [31:0] GEN_3760;
  reg [2:0] priority_44;
  reg [31:0] GEN_3761;
  reg [2:0] priority_45;
  reg [31:0] GEN_3762;
  reg [2:0] priority_46;
  reg [31:0] GEN_3763;
  reg [2:0] priority_47;
  reg [31:0] GEN_3764;
  reg [2:0] priority_48;
  reg [31:0] GEN_3765;
  reg [2:0] priority_49;
  reg [31:0] GEN_3766;
  reg [2:0] priority_50;
  reg [31:0] GEN_3767;
  reg [2:0] priority_51;
  reg [31:0] GEN_3768;
  reg [2:0] threshold_0;
  reg [31:0] GEN_3769;
  wire  T_2365_0;
  wire  T_2365_1;
  wire  T_2365_2;
  wire  T_2365_3;
  wire  T_2365_4;
  wire  T_2365_5;
  wire  T_2365_6;
  wire  T_2365_7;
  wire  T_2365_8;
  wire  T_2365_9;
  wire  T_2365_10;
  wire  T_2365_11;
  wire  T_2365_12;
  wire  T_2365_13;
  wire  T_2365_14;
  wire  T_2365_15;
  wire  T_2365_16;
  wire  T_2365_17;
  wire  T_2365_18;
  wire  T_2365_19;
  wire  T_2365_20;
  wire  T_2365_21;
  wire  T_2365_22;
  wire  T_2365_23;
  wire  T_2365_24;
  wire  T_2365_25;
  wire  T_2365_26;
  wire  T_2365_27;
  wire  T_2365_28;
  wire  T_2365_29;
  wire  T_2365_30;
  wire  T_2365_31;
  wire  T_2365_32;
  wire  T_2365_33;
  wire  T_2365_34;
  wire  T_2365_35;
  wire  T_2365_36;
  wire  T_2365_37;
  wire  T_2365_38;
  wire  T_2365_39;
  wire  T_2365_40;
  wire  T_2365_41;
  wire  T_2365_42;
  wire  T_2365_43;
  wire  T_2365_44;
  wire  T_2365_45;
  wire  T_2365_46;
  wire  T_2365_47;
  wire  T_2365_48;
  wire  T_2365_49;
  wire  T_2365_50;
  wire  T_2365_51;
  reg  pending_0;
  reg [31:0] GEN_3770;
  reg  pending_1;
  reg [31:0] GEN_3771;
  reg  pending_2;
  reg [31:0] GEN_3772;
  reg  pending_3;
  reg [31:0] GEN_3773;
  reg  pending_4;
  reg [31:0] GEN_3774;
  reg  pending_5;
  reg [31:0] GEN_3775;
  reg  pending_6;
  reg [31:0] GEN_3776;
  reg  pending_7;
  reg [31:0] GEN_3777;
  reg  pending_8;
  reg [31:0] GEN_3778;
  reg  pending_9;
  reg [31:0] GEN_3779;
  reg  pending_10;
  reg [31:0] GEN_3780;
  reg  pending_11;
  reg [31:0] GEN_3781;
  reg  pending_12;
  reg [31:0] GEN_3782;
  reg  pending_13;
  reg [31:0] GEN_3783;
  reg  pending_14;
  reg [31:0] GEN_3784;
  reg  pending_15;
  reg [31:0] GEN_3785;
  reg  pending_16;
  reg [31:0] GEN_3786;
  reg  pending_17;
  reg [31:0] GEN_3787;
  reg  pending_18;
  reg [31:0] GEN_3788;
  reg  pending_19;
  reg [31:0] GEN_3789;
  reg  pending_20;
  reg [31:0] GEN_3790;
  reg  pending_21;
  reg [31:0] GEN_3791;
  reg  pending_22;
  reg [31:0] GEN_3792;
  reg  pending_23;
  reg [31:0] GEN_3793;
  reg  pending_24;
  reg [31:0] GEN_3794;
  reg  pending_25;
  reg [31:0] GEN_3795;
  reg  pending_26;
  reg [31:0] GEN_3796;
  reg  pending_27;
  reg [31:0] GEN_3797;
  reg  pending_28;
  reg [31:0] GEN_3798;
  reg  pending_29;
  reg [31:0] GEN_3799;
  reg  pending_30;
  reg [31:0] GEN_3800;
  reg  pending_31;
  reg [31:0] GEN_3801;
  reg  pending_32;
  reg [31:0] GEN_3802;
  reg  pending_33;
  reg [31:0] GEN_3803;
  reg  pending_34;
  reg [31:0] GEN_3804;
  reg  pending_35;
  reg [31:0] GEN_3805;
  reg  pending_36;
  reg [31:0] GEN_3806;
  reg  pending_37;
  reg [31:0] GEN_3807;
  reg  pending_38;
  reg [31:0] GEN_3808;
  reg  pending_39;
  reg [31:0] GEN_3809;
  reg  pending_40;
  reg [31:0] GEN_3810;
  reg  pending_41;
  reg [31:0] GEN_3811;
  reg  pending_42;
  reg [31:0] GEN_3812;
  reg  pending_43;
  reg [31:0] GEN_3813;
  reg  pending_44;
  reg [31:0] GEN_3814;
  reg  pending_45;
  reg [31:0] GEN_3815;
  reg  pending_46;
  reg [31:0] GEN_3816;
  reg  pending_47;
  reg [31:0] GEN_3817;
  reg  pending_48;
  reg [31:0] GEN_3818;
  reg  pending_49;
  reg [31:0] GEN_3819;
  reg  pending_50;
  reg [31:0] GEN_3820;
  reg  pending_51;
  reg [31:0] GEN_3821;
  reg  enables_0_0;
  reg [31:0] GEN_3822;
  reg  enables_0_1;
  reg [31:0] GEN_3823;
  reg  enables_0_2;
  reg [31:0] GEN_3824;
  reg  enables_0_3;
  reg [31:0] GEN_3825;
  reg  enables_0_4;
  reg [31:0] GEN_3826;
  reg  enables_0_5;
  reg [31:0] GEN_3827;
  reg  enables_0_6;
  reg [31:0] GEN_3828;
  reg  enables_0_7;
  reg [31:0] GEN_3829;
  reg  enables_0_8;
  reg [31:0] GEN_3830;
  reg  enables_0_9;
  reg [31:0] GEN_3831;
  reg  enables_0_10;
  reg [31:0] GEN_3832;
  reg  enables_0_11;
  reg [31:0] GEN_3833;
  reg  enables_0_12;
  reg [31:0] GEN_3834;
  reg  enables_0_13;
  reg [31:0] GEN_3835;
  reg  enables_0_14;
  reg [31:0] GEN_3836;
  reg  enables_0_15;
  reg [31:0] GEN_3837;
  reg  enables_0_16;
  reg [31:0] GEN_3838;
  reg  enables_0_17;
  reg [31:0] GEN_3839;
  reg  enables_0_18;
  reg [31:0] GEN_3840;
  reg  enables_0_19;
  reg [31:0] GEN_3841;
  reg  enables_0_20;
  reg [31:0] GEN_3842;
  reg  enables_0_21;
  reg [31:0] GEN_3843;
  reg  enables_0_22;
  reg [31:0] GEN_3844;
  reg  enables_0_23;
  reg [31:0] GEN_3845;
  reg  enables_0_24;
  reg [31:0] GEN_3846;
  reg  enables_0_25;
  reg [31:0] GEN_3847;
  reg  enables_0_26;
  reg [31:0] GEN_3848;
  reg  enables_0_27;
  reg [31:0] GEN_3849;
  reg  enables_0_28;
  reg [31:0] GEN_3850;
  reg  enables_0_29;
  reg [31:0] GEN_3851;
  reg  enables_0_30;
  reg [31:0] GEN_3852;
  reg  enables_0_31;
  reg [31:0] GEN_3853;
  reg  enables_0_32;
  reg [31:0] GEN_3854;
  reg  enables_0_33;
  reg [31:0] GEN_3855;
  reg  enables_0_34;
  reg [31:0] GEN_3856;
  reg  enables_0_35;
  reg [31:0] GEN_3857;
  reg  enables_0_36;
  reg [31:0] GEN_3858;
  reg  enables_0_37;
  reg [31:0] GEN_3859;
  reg  enables_0_38;
  reg [31:0] GEN_3860;
  reg  enables_0_39;
  reg [31:0] GEN_3861;
  reg  enables_0_40;
  reg [31:0] GEN_3862;
  reg  enables_0_41;
  reg [31:0] GEN_3863;
  reg  enables_0_42;
  reg [31:0] GEN_3864;
  reg  enables_0_43;
  reg [31:0] GEN_3865;
  reg  enables_0_44;
  reg [31:0] GEN_3866;
  reg  enables_0_45;
  reg [31:0] GEN_3867;
  reg  enables_0_46;
  reg [31:0] GEN_3868;
  reg  enables_0_47;
  reg [31:0] GEN_3869;
  reg  enables_0_48;
  reg [31:0] GEN_3870;
  reg  enables_0_49;
  reg [31:0] GEN_3871;
  reg  enables_0_50;
  reg [31:0] GEN_3872;
  reg  enables_0_51;
  reg [31:0] GEN_3873;
  wire  T_2485;
  wire  GEN_9;
  wire  T_2489;
  wire  GEN_10;
  wire  T_2493;
  wire  GEN_11;
  wire  T_2497;
  wire  GEN_12;
  wire  T_2501;
  wire  GEN_13;
  wire  T_2505;
  wire  GEN_14;
  wire  T_2509;
  wire  GEN_15;
  wire  T_2513;
  wire  GEN_16;
  wire  T_2517;
  wire  GEN_17;
  wire  T_2521;
  wire  GEN_18;
  wire  T_2525;
  wire  GEN_19;
  wire  T_2529;
  wire  GEN_20;
  wire  T_2533;
  wire  GEN_21;
  wire  T_2537;
  wire  GEN_22;
  wire  T_2541;
  wire  GEN_23;
  wire  T_2545;
  wire  GEN_24;
  wire  T_2549;
  wire  GEN_25;
  wire  T_2553;
  wire  GEN_26;
  wire  T_2557;
  wire  GEN_27;
  wire  T_2561;
  wire  GEN_28;
  wire  T_2565;
  wire  GEN_29;
  wire  T_2569;
  wire  GEN_30;
  wire  T_2573;
  wire  GEN_31;
  wire  T_2577;
  wire  GEN_32;
  wire  T_2581;
  wire  GEN_33;
  wire  T_2585;
  wire  GEN_34;
  wire  T_2589;
  wire  GEN_35;
  wire  T_2593;
  wire  GEN_36;
  wire  T_2597;
  wire  GEN_37;
  wire  T_2601;
  wire  GEN_38;
  wire  T_2605;
  wire  GEN_39;
  wire  T_2609;
  wire  GEN_40;
  wire  T_2613;
  wire  GEN_41;
  wire  T_2617;
  wire  GEN_42;
  wire  T_2621;
  wire  GEN_43;
  wire  T_2625;
  wire  GEN_44;
  wire  T_2629;
  wire  GEN_45;
  wire  T_2633;
  wire  GEN_46;
  wire  T_2637;
  wire  GEN_47;
  wire  T_2641;
  wire  GEN_48;
  wire  T_2645;
  wire  GEN_49;
  wire  T_2649;
  wire  GEN_50;
  wire  T_2653;
  wire  GEN_51;
  wire  T_2657;
  wire  GEN_52;
  wire  T_2661;
  wire  GEN_53;
  wire  T_2665;
  wire  GEN_54;
  wire  T_2669;
  wire  GEN_55;
  wire  T_2673;
  wire  GEN_56;
  wire  T_2677;
  wire  GEN_57;
  wire  T_2681;
  wire  GEN_58;
  wire  T_2685;
  wire  GEN_59;
  reg [5:0] maxDevs_0;
  reg [31:0] GEN_3874;
  wire  T_2692;
  wire [3:0] T_2693;
  wire  T_2694;
  wire [3:0] T_2695;
  wire  T_2696;
  wire [3:0] T_2697;
  wire  T_2698;
  wire [3:0] T_2699;
  wire  T_2700;
  wire [3:0] T_2701;
  wire  T_2702;
  wire [3:0] T_2703;
  wire  T_2704;
  wire [3:0] T_2705;
  wire  T_2706;
  wire [3:0] T_2707;
  wire  T_2708;
  wire [3:0] T_2709;
  wire  T_2710;
  wire [3:0] T_2711;
  wire  T_2712;
  wire [3:0] T_2713;
  wire  T_2714;
  wire [3:0] T_2715;
  wire  T_2716;
  wire [3:0] T_2717;
  wire  T_2718;
  wire [3:0] T_2719;
  wire  T_2720;
  wire [3:0] T_2721;
  wire  T_2722;
  wire [3:0] T_2723;
  wire  T_2724;
  wire [3:0] T_2725;
  wire  T_2726;
  wire [3:0] T_2727;
  wire  T_2728;
  wire [3:0] T_2729;
  wire  T_2730;
  wire [3:0] T_2731;
  wire  T_2732;
  wire [3:0] T_2733;
  wire  T_2734;
  wire [3:0] T_2735;
  wire  T_2736;
  wire [3:0] T_2737;
  wire  T_2738;
  wire [3:0] T_2739;
  wire  T_2740;
  wire [3:0] T_2741;
  wire  T_2742;
  wire [3:0] T_2743;
  wire  T_2744;
  wire [3:0] T_2745;
  wire  T_2746;
  wire [3:0] T_2747;
  wire  T_2748;
  wire [3:0] T_2749;
  wire  T_2750;
  wire [3:0] T_2751;
  wire  T_2752;
  wire [3:0] T_2753;
  wire  T_2754;
  wire [3:0] T_2755;
  wire  T_2756;
  wire [3:0] T_2757;
  wire  T_2758;
  wire [3:0] T_2759;
  wire  T_2760;
  wire [3:0] T_2761;
  wire  T_2762;
  wire [3:0] T_2763;
  wire  T_2764;
  wire [3:0] T_2765;
  wire  T_2766;
  wire [3:0] T_2767;
  wire  T_2768;
  wire [3:0] T_2769;
  wire  T_2770;
  wire [3:0] T_2771;
  wire  T_2772;
  wire [3:0] T_2773;
  wire  T_2774;
  wire [3:0] T_2775;
  wire  T_2776;
  wire [3:0] T_2777;
  wire  T_2778;
  wire [3:0] T_2779;
  wire  T_2780;
  wire [3:0] T_2781;
  wire  T_2782;
  wire [3:0] T_2783;
  wire  T_2784;
  wire [3:0] T_2785;
  wire  T_2786;
  wire [3:0] T_2787;
  wire  T_2788;
  wire [3:0] T_2789;
  wire  T_2790;
  wire [3:0] T_2791;
  wire  T_2792;
  wire [3:0] T_2793;
  wire  T_2798;
  wire [3:0] T_2799;
  wire  T_2802;
  wire  T_2805;
  wire [3:0] T_2806;
  wire  T_2809;
  wire  T_2810;
  wire [3:0] T_2811;
  wire [1:0] GEN_3489;
  wire [1:0] T_2813;
  wire [1:0] T_2814;
  wire  T_2817;
  wire [3:0] T_2818;
  wire  T_2821;
  wire  T_2824;
  wire [3:0] T_2825;
  wire  T_2828;
  wire  T_2829;
  wire [3:0] T_2830;
  wire [1:0] GEN_3490;
  wire [1:0] T_2832;
  wire [1:0] T_2833;
  wire  T_2834;
  wire [3:0] T_2835;
  wire [2:0] GEN_3491;
  wire [2:0] T_2837;
  wire [2:0] T_2838;
  wire  T_2841;
  wire [3:0] T_2842;
  wire  T_2845;
  wire  T_2848;
  wire [3:0] T_2849;
  wire  T_2852;
  wire  T_2853;
  wire [3:0] T_2854;
  wire [1:0] GEN_3492;
  wire [1:0] T_2856;
  wire [1:0] T_2857;
  wire  T_2860;
  wire [3:0] T_2861;
  wire  T_2864;
  wire  T_2867;
  wire [3:0] T_2868;
  wire  T_2871;
  wire  T_2872;
  wire [3:0] T_2873;
  wire [1:0] GEN_3493;
  wire [1:0] T_2875;
  wire [1:0] T_2876;
  wire  T_2877;
  wire [3:0] T_2878;
  wire [2:0] GEN_3494;
  wire [2:0] T_2880;
  wire [2:0] T_2881;
  wire  T_2882;
  wire [3:0] T_2883;
  wire [3:0] GEN_3495;
  wire [3:0] T_2885;
  wire [3:0] T_2886;
  wire  T_2889;
  wire [3:0] T_2890;
  wire  T_2893;
  wire  T_2896;
  wire [3:0] T_2897;
  wire  T_2900;
  wire  T_2901;
  wire [3:0] T_2902;
  wire [1:0] GEN_3496;
  wire [1:0] T_2904;
  wire [1:0] T_2905;
  wire  T_2908;
  wire [3:0] T_2909;
  wire  T_2912;
  wire  T_2915;
  wire [3:0] T_2916;
  wire  T_2919;
  wire  T_2920;
  wire [3:0] T_2921;
  wire [1:0] GEN_3497;
  wire [1:0] T_2923;
  wire [1:0] T_2924;
  wire  T_2925;
  wire [3:0] T_2926;
  wire [2:0] GEN_3498;
  wire [2:0] T_2928;
  wire [2:0] T_2929;
  wire  T_2932;
  wire [3:0] T_2933;
  wire  T_2936;
  wire  T_2939;
  wire [3:0] T_2940;
  wire  T_2943;
  wire  T_2944;
  wire [3:0] T_2945;
  wire [1:0] GEN_3499;
  wire [1:0] T_2947;
  wire [1:0] T_2948;
  wire  T_2951;
  wire [3:0] T_2952;
  wire  T_2955;
  wire  T_2958;
  wire [3:0] T_2959;
  wire  T_2962;
  wire  T_2963;
  wire [3:0] T_2964;
  wire [1:0] GEN_3500;
  wire [1:0] T_2966;
  wire [1:0] T_2967;
  wire  T_2968;
  wire [3:0] T_2969;
  wire [2:0] GEN_3501;
  wire [2:0] T_2971;
  wire [2:0] T_2972;
  wire  T_2973;
  wire [3:0] T_2974;
  wire [3:0] GEN_3502;
  wire [3:0] T_2976;
  wire [3:0] T_2977;
  wire  T_2978;
  wire [3:0] T_2979;
  wire [4:0] GEN_3503;
  wire [4:0] T_2981;
  wire [4:0] T_2982;
  wire  T_2985;
  wire [3:0] T_2986;
  wire  T_2989;
  wire  T_2992;
  wire [3:0] T_2993;
  wire  T_2996;
  wire  T_2997;
  wire [3:0] T_2998;
  wire [1:0] GEN_3504;
  wire [1:0] T_3000;
  wire [1:0] T_3001;
  wire  T_3004;
  wire [3:0] T_3005;
  wire  T_3008;
  wire  T_3011;
  wire [3:0] T_3012;
  wire  T_3015;
  wire  T_3016;
  wire [3:0] T_3017;
  wire [1:0] GEN_3505;
  wire [1:0] T_3019;
  wire [1:0] T_3020;
  wire  T_3021;
  wire [3:0] T_3022;
  wire [2:0] GEN_3506;
  wire [2:0] T_3024;
  wire [2:0] T_3025;
  wire  T_3028;
  wire [3:0] T_3029;
  wire  T_3032;
  wire  T_3035;
  wire [3:0] T_3036;
  wire  T_3039;
  wire  T_3040;
  wire [3:0] T_3041;
  wire [1:0] GEN_3507;
  wire [1:0] T_3043;
  wire [1:0] T_3044;
  wire  T_3047;
  wire [3:0] T_3048;
  wire  T_3051;
  wire  T_3054;
  wire [3:0] T_3055;
  wire  T_3058;
  wire  T_3059;
  wire [3:0] T_3060;
  wire [1:0] GEN_3508;
  wire [1:0] T_3062;
  wire [1:0] T_3063;
  wire  T_3064;
  wire [3:0] T_3065;
  wire [2:0] GEN_3509;
  wire [2:0] T_3067;
  wire [2:0] T_3068;
  wire  T_3069;
  wire [3:0] T_3070;
  wire [3:0] GEN_3510;
  wire [3:0] T_3072;
  wire [3:0] T_3073;
  wire  T_3076;
  wire [3:0] T_3077;
  wire  T_3080;
  wire  T_3083;
  wire [3:0] T_3084;
  wire  T_3087;
  wire  T_3088;
  wire [3:0] T_3089;
  wire [1:0] GEN_3511;
  wire [1:0] T_3091;
  wire [1:0] T_3092;
  wire  T_3093;
  wire [3:0] T_3094;
  wire [4:0] GEN_3512;
  wire [4:0] T_3096;
  wire [4:0] T_3097;
  wire  T_3098;
  wire [3:0] T_3099;
  wire [5:0] GEN_3513;
  wire [5:0] T_3101;
  wire [5:0] T_3102;
  reg [3:0] T_3103;
  reg [31:0] GEN_3875;
  wire [3:0] T_3105;
  wire  T_3106;
  wire  T_3130_ready;
  wire  T_3130_valid;
  wire  T_3130_bits_read;
  wire [23:0] T_3130_bits_index;
  wire [31:0] T_3130_bits_data;
  wire [3:0] T_3130_bits_mask;
  wire [9:0] T_3130_bits_extra;
  wire  T_3147;
  wire [25:0] T_3148;
  wire [1:0] T_3149;
  wire [6:0] T_3150;
  wire [9:0] T_3151;
  wire  T_3169_ready;
  wire  T_3169_valid;
  wire  T_3169_bits_read;
  wire [31:0] T_3169_bits_data;
  wire [9:0] T_3169_bits_extra;
  wire  T_3205_ready;
  wire  T_3205_valid;
  wire  T_3205_bits_read;
  wire [23:0] T_3205_bits_index;
  wire [31:0] T_3205_bits_data;
  wire [3:0] T_3205_bits_mask;
  wire [9:0] T_3205_bits_extra;
  wire  T_4309_0;
  wire  T_4309_1;
  wire  T_4309_2;
  wire  T_4309_3;
  wire  T_4309_4;
  wire  T_4309_5;
  wire  T_4309_6;
  wire  T_4309_7;
  wire  T_4309_8;
  wire  T_4309_9;
  wire  T_4309_10;
  wire  T_4309_11;
  wire  T_4309_12;
  wire  T_4309_13;
  wire  T_4309_14;
  wire  T_4309_15;
  wire  T_4309_16;
  wire  T_4309_17;
  wire  T_4309_18;
  wire  T_4309_19;
  wire  T_4309_20;
  wire  T_4309_21;
  wire  T_4309_22;
  wire  T_4309_23;
  wire  T_4309_24;
  wire  T_4309_25;
  wire  T_4309_26;
  wire  T_4309_27;
  wire  T_4309_28;
  wire  T_4309_29;
  wire  T_4309_30;
  wire  T_4309_31;
  wire  T_4309_32;
  wire  T_4309_33;
  wire  T_4309_34;
  wire  T_4309_35;
  wire  T_4309_36;
  wire  T_4309_37;
  wire  T_4309_38;
  wire  T_4309_39;
  wire  T_4309_40;
  wire  T_4309_41;
  wire  T_4309_42;
  wire  T_4309_43;
  wire  T_4309_44;
  wire  T_4309_45;
  wire  T_4309_46;
  wire  T_4309_47;
  wire  T_4309_48;
  wire  T_4309_49;
  wire  T_4309_50;
  wire  T_4309_51;
  wire  T_4309_52;
  wire  T_4309_53;
  wire  T_4309_54;
  wire  T_4309_55;
  wire  T_4309_56;
  wire  T_4309_57;
  wire  T_4309_58;
  wire  T_4309_59;
  wire  T_4309_60;
  wire  T_4309_61;
  wire  T_4309_62;
  wire  T_4309_63;
  wire  T_4309_64;
  wire  T_4309_65;
  wire  T_4309_66;
  wire  T_4309_67;
  wire  T_4309_68;
  wire  T_4309_69;
  wire  T_4309_70;
  wire  T_4309_71;
  wire  T_4309_72;
  wire  T_4309_73;
  wire  T_4309_74;
  wire  T_4309_75;
  wire  T_4309_76;
  wire  T_4309_77;
  wire  T_4309_78;
  wire  T_4309_79;
  wire  T_4309_80;
  wire  T_4309_81;
  wire  T_4309_82;
  wire  T_4309_83;
  wire  T_4309_84;
  wire  T_4309_85;
  wire  T_4309_86;
  wire  T_4309_87;
  wire  T_4309_88;
  wire  T_4309_89;
  wire  T_4309_90;
  wire  T_4309_91;
  wire  T_4309_92;
  wire  T_4309_93;
  wire  T_4309_94;
  wire  T_4309_95;
  wire  T_4309_96;
  wire  T_4309_97;
  wire  T_4309_98;
  wire  T_4309_99;
  wire  T_4309_100;
  wire  T_4309_101;
  wire  T_4309_102;
  wire  T_4309_103;
  wire  T_4309_104;
  wire  T_4309_105;
  wire  T_4309_106;
  wire  T_4309_107;
  wire  T_4309_108;
  wire  T_4309_109;
  wire  T_4309_110;
  wire  T_4309_111;
  wire  T_4309_112;
  wire  T_4309_113;
  wire  T_4309_114;
  wire  T_4309_115;
  wire  T_4309_116;
  wire  T_4309_117;
  wire  T_4309_118;
  wire  T_4309_119;
  wire  T_4309_120;
  wire  T_4309_121;
  wire  T_4309_122;
  wire  T_4309_123;
  wire  T_4309_124;
  wire  T_4309_125;
  wire  T_4309_126;
  wire  T_4309_127;
  wire  T_4309_128;
  wire  T_4309_129;
  wire  T_4309_130;
  wire  T_4309_131;
  wire  T_4309_132;
  wire  T_4309_133;
  wire  T_4309_134;
  wire  T_4309_135;
  wire  T_4309_136;
  wire  T_4309_137;
  wire  T_4309_138;
  wire  T_4309_139;
  wire  T_4309_140;
  wire  T_4309_141;
  wire  T_4309_142;
  wire  T_4309_143;
  wire  T_4309_144;
  wire  T_4309_145;
  wire  T_4309_146;
  wire  T_4309_147;
  wire  T_4309_148;
  wire  T_4309_149;
  wire  T_4309_150;
  wire  T_4309_151;
  wire  T_4309_152;
  wire  T_4309_153;
  wire  T_4309_154;
  wire  T_4309_155;
  wire  T_4309_156;
  wire  T_4309_157;
  wire  T_4314_0;
  wire  T_4314_1;
  wire  T_4314_2;
  wire  T_4314_3;
  wire  T_4314_4;
  wire  T_4314_5;
  wire  T_4314_6;
  wire  T_4314_7;
  wire  T_4314_8;
  wire  T_4314_9;
  wire  T_4314_10;
  wire  T_4314_11;
  wire  T_4314_12;
  wire  T_4314_13;
  wire  T_4314_14;
  wire  T_4314_15;
  wire  T_4314_16;
  wire  T_4314_17;
  wire  T_4314_18;
  wire  T_4314_19;
  wire  T_4314_20;
  wire  T_4314_21;
  wire  T_4314_22;
  wire  T_4314_23;
  wire  T_4314_24;
  wire  T_4314_25;
  wire  T_4314_26;
  wire  T_4314_27;
  wire  T_4314_28;
  wire  T_4314_29;
  wire  T_4314_30;
  wire  T_4314_31;
  wire  T_4314_32;
  wire  T_4314_33;
  wire  T_4314_34;
  wire  T_4314_35;
  wire  T_4314_36;
  wire  T_4314_37;
  wire  T_4314_38;
  wire  T_4314_39;
  wire  T_4314_40;
  wire  T_4314_41;
  wire  T_4314_42;
  wire  T_4314_43;
  wire  T_4314_44;
  wire  T_4314_45;
  wire  T_4314_46;
  wire  T_4314_47;
  wire  T_4314_48;
  wire  T_4314_49;
  wire  T_4314_50;
  wire  T_4314_51;
  wire  T_4314_52;
  wire  T_4314_53;
  wire  T_4314_54;
  wire  T_4314_55;
  wire  T_4314_56;
  wire  T_4314_57;
  wire  T_4314_58;
  wire  T_4314_59;
  wire  T_4314_60;
  wire  T_4314_61;
  wire  T_4314_62;
  wire  T_4314_63;
  wire  T_4314_64;
  wire  T_4314_65;
  wire  T_4314_66;
  wire  T_4314_67;
  wire  T_4314_68;
  wire  T_4314_69;
  wire  T_4314_70;
  wire  T_4314_71;
  wire  T_4314_72;
  wire  T_4314_73;
  wire  T_4314_74;
  wire  T_4314_75;
  wire  T_4314_76;
  wire  T_4314_77;
  wire  T_4314_78;
  wire  T_4314_79;
  wire  T_4314_80;
  wire  T_4314_81;
  wire  T_4314_82;
  wire  T_4314_83;
  wire  T_4314_84;
  wire  T_4314_85;
  wire  T_4314_86;
  wire  T_4314_87;
  wire  T_4314_88;
  wire  T_4314_89;
  wire  T_4314_90;
  wire  T_4314_91;
  wire  T_4314_92;
  wire  T_4314_93;
  wire  T_4314_94;
  wire  T_4314_95;
  wire  T_4314_96;
  wire  T_4314_97;
  wire  T_4314_98;
  wire  T_4314_99;
  wire  T_4314_100;
  wire  T_4314_101;
  wire  T_4314_102;
  wire  T_4314_103;
  wire  T_4314_104;
  wire  T_4314_105;
  wire  T_4314_106;
  wire  T_4314_107;
  wire  T_4314_108;
  wire  T_4314_109;
  wire  T_4314_110;
  wire  T_4314_111;
  wire  T_4314_112;
  wire  T_4314_113;
  wire  T_4314_114;
  wire  T_4314_115;
  wire  T_4314_116;
  wire  T_4314_117;
  wire  T_4314_118;
  wire  T_4314_119;
  wire  T_4314_120;
  wire  T_4314_121;
  wire  T_4314_122;
  wire  T_4314_123;
  wire  T_4314_124;
  wire  T_4314_125;
  wire  T_4314_126;
  wire  T_4314_127;
  wire  T_4314_128;
  wire  T_4314_129;
  wire  T_4314_130;
  wire  T_4314_131;
  wire  T_4314_132;
  wire  T_4314_133;
  wire  T_4314_134;
  wire  T_4314_135;
  wire  T_4314_136;
  wire  T_4314_137;
  wire  T_4314_138;
  wire  T_4314_139;
  wire  T_4314_140;
  wire  T_4314_141;
  wire  T_4314_142;
  wire  T_4314_143;
  wire  T_4314_144;
  wire  T_4314_145;
  wire  T_4314_146;
  wire  T_4314_147;
  wire  T_4314_148;
  wire  T_4314_149;
  wire  T_4314_150;
  wire  T_4314_151;
  wire  T_4314_152;
  wire  T_4314_153;
  wire  T_4314_154;
  wire  T_4314_155;
  wire  T_4314_156;
  wire  T_4314_157;
  wire  T_4319_0;
  wire  T_4319_1;
  wire  T_4319_2;
  wire  T_4319_3;
  wire  T_4319_4;
  wire  T_4319_5;
  wire  T_4319_6;
  wire  T_4319_7;
  wire  T_4319_8;
  wire  T_4319_9;
  wire  T_4319_10;
  wire  T_4319_11;
  wire  T_4319_12;
  wire  T_4319_13;
  wire  T_4319_14;
  wire  T_4319_15;
  wire  T_4319_16;
  wire  T_4319_17;
  wire  T_4319_18;
  wire  T_4319_19;
  wire  T_4319_20;
  wire  T_4319_21;
  wire  T_4319_22;
  wire  T_4319_23;
  wire  T_4319_24;
  wire  T_4319_25;
  wire  T_4319_26;
  wire  T_4319_27;
  wire  T_4319_28;
  wire  T_4319_29;
  wire  T_4319_30;
  wire  T_4319_31;
  wire  T_4319_32;
  wire  T_4319_33;
  wire  T_4319_34;
  wire  T_4319_35;
  wire  T_4319_36;
  wire  T_4319_37;
  wire  T_4319_38;
  wire  T_4319_39;
  wire  T_4319_40;
  wire  T_4319_41;
  wire  T_4319_42;
  wire  T_4319_43;
  wire  T_4319_44;
  wire  T_4319_45;
  wire  T_4319_46;
  wire  T_4319_47;
  wire  T_4319_48;
  wire  T_4319_49;
  wire  T_4319_50;
  wire  T_4319_51;
  wire  T_4319_52;
  wire  T_4319_53;
  wire  T_4319_54;
  wire  T_4319_55;
  wire  T_4319_56;
  wire  T_4319_57;
  wire  T_4319_58;
  wire  T_4319_59;
  wire  T_4319_60;
  wire  T_4319_61;
  wire  T_4319_62;
  wire  T_4319_63;
  wire  T_4319_64;
  wire  T_4319_65;
  wire  T_4319_66;
  wire  T_4319_67;
  wire  T_4319_68;
  wire  T_4319_69;
  wire  T_4319_70;
  wire  T_4319_71;
  wire  T_4319_72;
  wire  T_4319_73;
  wire  T_4319_74;
  wire  T_4319_75;
  wire  T_4319_76;
  wire  T_4319_77;
  wire  T_4319_78;
  wire  T_4319_79;
  wire  T_4319_80;
  wire  T_4319_81;
  wire  T_4319_82;
  wire  T_4319_83;
  wire  T_4319_84;
  wire  T_4319_85;
  wire  T_4319_86;
  wire  T_4319_87;
  wire  T_4319_88;
  wire  T_4319_89;
  wire  T_4319_90;
  wire  T_4319_91;
  wire  T_4319_92;
  wire  T_4319_93;
  wire  T_4319_94;
  wire  T_4319_95;
  wire  T_4319_96;
  wire  T_4319_97;
  wire  T_4319_98;
  wire  T_4319_99;
  wire  T_4319_100;
  wire  T_4319_101;
  wire  T_4319_102;
  wire  T_4319_103;
  wire  T_4319_104;
  wire  T_4319_105;
  wire  T_4319_106;
  wire  T_4319_107;
  wire  T_4319_108;
  wire  T_4319_109;
  wire  T_4319_110;
  wire  T_4319_111;
  wire  T_4319_112;
  wire  T_4319_113;
  wire  T_4319_114;
  wire  T_4319_115;
  wire  T_4319_116;
  wire  T_4319_117;
  wire  T_4319_118;
  wire  T_4319_119;
  wire  T_4319_120;
  wire  T_4319_121;
  wire  T_4319_122;
  wire  T_4319_123;
  wire  T_4319_124;
  wire  T_4319_125;
  wire  T_4319_126;
  wire  T_4319_127;
  wire  T_4319_128;
  wire  T_4319_129;
  wire  T_4319_130;
  wire  T_4319_131;
  wire  T_4319_132;
  wire  T_4319_133;
  wire  T_4319_134;
  wire  T_4319_135;
  wire  T_4319_136;
  wire  T_4319_137;
  wire  T_4319_138;
  wire  T_4319_139;
  wire  T_4319_140;
  wire  T_4319_141;
  wire  T_4319_142;
  wire  T_4319_143;
  wire  T_4319_144;
  wire  T_4319_145;
  wire  T_4319_146;
  wire  T_4319_147;
  wire  T_4319_148;
  wire  T_4319_149;
  wire  T_4319_150;
  wire  T_4319_151;
  wire  T_4319_152;
  wire  T_4319_153;
  wire  T_4319_154;
  wire  T_4319_155;
  wire  T_4319_156;
  wire  T_4319_157;
  wire  T_4324_0;
  wire  T_4324_1;
  wire  T_4324_2;
  wire  T_4324_3;
  wire  T_4324_4;
  wire  T_4324_5;
  wire  T_4324_6;
  wire  T_4324_7;
  wire  T_4324_8;
  wire  T_4324_9;
  wire  T_4324_10;
  wire  T_4324_11;
  wire  T_4324_12;
  wire  T_4324_13;
  wire  T_4324_14;
  wire  T_4324_15;
  wire  T_4324_16;
  wire  T_4324_17;
  wire  T_4324_18;
  wire  T_4324_19;
  wire  T_4324_20;
  wire  T_4324_21;
  wire  T_4324_22;
  wire  T_4324_23;
  wire  T_4324_24;
  wire  T_4324_25;
  wire  T_4324_26;
  wire  T_4324_27;
  wire  T_4324_28;
  wire  T_4324_29;
  wire  T_4324_30;
  wire  T_4324_31;
  wire  T_4324_32;
  wire  T_4324_33;
  wire  T_4324_34;
  wire  T_4324_35;
  wire  T_4324_36;
  wire  T_4324_37;
  wire  T_4324_38;
  wire  T_4324_39;
  wire  T_4324_40;
  wire  T_4324_41;
  wire  T_4324_42;
  wire  T_4324_43;
  wire  T_4324_44;
  wire  T_4324_45;
  wire  T_4324_46;
  wire  T_4324_47;
  wire  T_4324_48;
  wire  T_4324_49;
  wire  T_4324_50;
  wire  T_4324_51;
  wire  T_4324_52;
  wire  T_4324_53;
  wire  T_4324_54;
  wire  T_4324_55;
  wire  T_4324_56;
  wire  T_4324_57;
  wire  T_4324_58;
  wire  T_4324_59;
  wire  T_4324_60;
  wire  T_4324_61;
  wire  T_4324_62;
  wire  T_4324_63;
  wire  T_4324_64;
  wire  T_4324_65;
  wire  T_4324_66;
  wire  T_4324_67;
  wire  T_4324_68;
  wire  T_4324_69;
  wire  T_4324_70;
  wire  T_4324_71;
  wire  T_4324_72;
  wire  T_4324_73;
  wire  T_4324_74;
  wire  T_4324_75;
  wire  T_4324_76;
  wire  T_4324_77;
  wire  T_4324_78;
  wire  T_4324_79;
  wire  T_4324_80;
  wire  T_4324_81;
  wire  T_4324_82;
  wire  T_4324_83;
  wire  T_4324_84;
  wire  T_4324_85;
  wire  T_4324_86;
  wire  T_4324_87;
  wire  T_4324_88;
  wire  T_4324_89;
  wire  T_4324_90;
  wire  T_4324_91;
  wire  T_4324_92;
  wire  T_4324_93;
  wire  T_4324_94;
  wire  T_4324_95;
  wire  T_4324_96;
  wire  T_4324_97;
  wire  T_4324_98;
  wire  T_4324_99;
  wire  T_4324_100;
  wire  T_4324_101;
  wire  T_4324_102;
  wire  T_4324_103;
  wire  T_4324_104;
  wire  T_4324_105;
  wire  T_4324_106;
  wire  T_4324_107;
  wire  T_4324_108;
  wire  T_4324_109;
  wire  T_4324_110;
  wire  T_4324_111;
  wire  T_4324_112;
  wire  T_4324_113;
  wire  T_4324_114;
  wire  T_4324_115;
  wire  T_4324_116;
  wire  T_4324_117;
  wire  T_4324_118;
  wire  T_4324_119;
  wire  T_4324_120;
  wire  T_4324_121;
  wire  T_4324_122;
  wire  T_4324_123;
  wire  T_4324_124;
  wire  T_4324_125;
  wire  T_4324_126;
  wire  T_4324_127;
  wire  T_4324_128;
  wire  T_4324_129;
  wire  T_4324_130;
  wire  T_4324_131;
  wire  T_4324_132;
  wire  T_4324_133;
  wire  T_4324_134;
  wire  T_4324_135;
  wire  T_4324_136;
  wire  T_4324_137;
  wire  T_4324_138;
  wire  T_4324_139;
  wire  T_4324_140;
  wire  T_4324_141;
  wire  T_4324_142;
  wire  T_4324_143;
  wire  T_4324_144;
  wire  T_4324_145;
  wire  T_4324_146;
  wire  T_4324_147;
  wire  T_4324_148;
  wire  T_4324_149;
  wire  T_4324_150;
  wire  T_4324_151;
  wire  T_4324_152;
  wire  T_4324_153;
  wire  T_4324_154;
  wire  T_4324_155;
  wire  T_4324_156;
  wire  T_4324_157;
  wire  T_4329_0;
  wire  T_4329_1;
  wire  T_4329_2;
  wire  T_4329_3;
  wire  T_4329_4;
  wire  T_4329_5;
  wire  T_4329_6;
  wire  T_4329_7;
  wire  T_4329_8;
  wire  T_4329_9;
  wire  T_4329_10;
  wire  T_4329_11;
  wire  T_4329_12;
  wire  T_4329_13;
  wire  T_4329_14;
  wire  T_4329_15;
  wire  T_4329_16;
  wire  T_4329_17;
  wire  T_4329_18;
  wire  T_4329_19;
  wire  T_4329_20;
  wire  T_4329_21;
  wire  T_4329_22;
  wire  T_4329_23;
  wire  T_4329_24;
  wire  T_4329_25;
  wire  T_4329_26;
  wire  T_4329_27;
  wire  T_4329_28;
  wire  T_4329_29;
  wire  T_4329_30;
  wire  T_4329_31;
  wire  T_4329_32;
  wire  T_4329_33;
  wire  T_4329_34;
  wire  T_4329_35;
  wire  T_4329_36;
  wire  T_4329_37;
  wire  T_4329_38;
  wire  T_4329_39;
  wire  T_4329_40;
  wire  T_4329_41;
  wire  T_4329_42;
  wire  T_4329_43;
  wire  T_4329_44;
  wire  T_4329_45;
  wire  T_4329_46;
  wire  T_4329_47;
  wire  T_4329_48;
  wire  T_4329_49;
  wire  T_4329_50;
  wire  T_4329_51;
  wire  T_4329_52;
  wire  T_4329_53;
  wire  T_4329_54;
  wire  T_4329_55;
  wire  T_4329_56;
  wire  T_4329_57;
  wire  T_4329_58;
  wire  T_4329_59;
  wire  T_4329_60;
  wire  T_4329_61;
  wire  T_4329_62;
  wire  T_4329_63;
  wire  T_4329_64;
  wire  T_4329_65;
  wire  T_4329_66;
  wire  T_4329_67;
  wire  T_4329_68;
  wire  T_4329_69;
  wire  T_4329_70;
  wire  T_4329_71;
  wire  T_4329_72;
  wire  T_4329_73;
  wire  T_4329_74;
  wire  T_4329_75;
  wire  T_4329_76;
  wire  T_4329_77;
  wire  T_4329_78;
  wire  T_4329_79;
  wire  T_4329_80;
  wire  T_4329_81;
  wire  T_4329_82;
  wire  T_4329_83;
  wire  T_4329_84;
  wire  T_4329_85;
  wire  T_4329_86;
  wire  T_4329_87;
  wire  T_4329_88;
  wire  T_4329_89;
  wire  T_4329_90;
  wire  T_4329_91;
  wire  T_4329_92;
  wire  T_4329_93;
  wire  T_4329_94;
  wire  T_4329_95;
  wire  T_4329_96;
  wire  T_4329_97;
  wire  T_4329_98;
  wire  T_4329_99;
  wire  T_4329_100;
  wire  T_4329_101;
  wire  T_4329_102;
  wire  T_4329_103;
  wire  T_4329_104;
  wire  T_4329_105;
  wire  T_4329_106;
  wire  T_4329_107;
  wire  T_4329_108;
  wire  T_4329_109;
  wire  T_4329_110;
  wire  T_4329_111;
  wire  T_4329_112;
  wire  T_4329_113;
  wire  T_4329_114;
  wire  T_4329_115;
  wire  T_4329_116;
  wire  T_4329_117;
  wire  T_4329_118;
  wire  T_4329_119;
  wire  T_4329_120;
  wire  T_4329_121;
  wire  T_4329_122;
  wire  T_4329_123;
  wire  T_4329_124;
  wire  T_4329_125;
  wire  T_4329_126;
  wire  T_4329_127;
  wire  T_4329_128;
  wire  T_4329_129;
  wire  T_4329_130;
  wire  T_4329_131;
  wire  T_4329_132;
  wire  T_4329_133;
  wire  T_4329_134;
  wire  T_4329_135;
  wire  T_4329_136;
  wire  T_4329_137;
  wire  T_4329_138;
  wire  T_4329_139;
  wire  T_4329_140;
  wire  T_4329_141;
  wire  T_4329_142;
  wire  T_4329_143;
  wire  T_4329_144;
  wire  T_4329_145;
  wire  T_4329_146;
  wire  T_4329_147;
  wire  T_4329_148;
  wire  T_4329_149;
  wire  T_4329_150;
  wire  T_4329_151;
  wire  T_4329_152;
  wire  T_4329_153;
  wire  T_4329_154;
  wire  T_4329_155;
  wire  T_4329_156;
  wire  T_4329_157;
  wire  T_4334_0;
  wire  T_4334_1;
  wire  T_4334_2;
  wire  T_4334_3;
  wire  T_4334_4;
  wire  T_4334_5;
  wire  T_4334_6;
  wire  T_4334_7;
  wire  T_4334_8;
  wire  T_4334_9;
  wire  T_4334_10;
  wire  T_4334_11;
  wire  T_4334_12;
  wire  T_4334_13;
  wire  T_4334_14;
  wire  T_4334_15;
  wire  T_4334_16;
  wire  T_4334_17;
  wire  T_4334_18;
  wire  T_4334_19;
  wire  T_4334_20;
  wire  T_4334_21;
  wire  T_4334_22;
  wire  T_4334_23;
  wire  T_4334_24;
  wire  T_4334_25;
  wire  T_4334_26;
  wire  T_4334_27;
  wire  T_4334_28;
  wire  T_4334_29;
  wire  T_4334_30;
  wire  T_4334_31;
  wire  T_4334_32;
  wire  T_4334_33;
  wire  T_4334_34;
  wire  T_4334_35;
  wire  T_4334_36;
  wire  T_4334_37;
  wire  T_4334_38;
  wire  T_4334_39;
  wire  T_4334_40;
  wire  T_4334_41;
  wire  T_4334_42;
  wire  T_4334_43;
  wire  T_4334_44;
  wire  T_4334_45;
  wire  T_4334_46;
  wire  T_4334_47;
  wire  T_4334_48;
  wire  T_4334_49;
  wire  T_4334_50;
  wire  T_4334_51;
  wire  T_4334_52;
  wire  T_4334_53;
  wire  T_4334_54;
  wire  T_4334_55;
  wire  T_4334_56;
  wire  T_4334_57;
  wire  T_4334_58;
  wire  T_4334_59;
  wire  T_4334_60;
  wire  T_4334_61;
  wire  T_4334_62;
  wire  T_4334_63;
  wire  T_4334_64;
  wire  T_4334_65;
  wire  T_4334_66;
  wire  T_4334_67;
  wire  T_4334_68;
  wire  T_4334_69;
  wire  T_4334_70;
  wire  T_4334_71;
  wire  T_4334_72;
  wire  T_4334_73;
  wire  T_4334_74;
  wire  T_4334_75;
  wire  T_4334_76;
  wire  T_4334_77;
  wire  T_4334_78;
  wire  T_4334_79;
  wire  T_4334_80;
  wire  T_4334_81;
  wire  T_4334_82;
  wire  T_4334_83;
  wire  T_4334_84;
  wire  T_4334_85;
  wire  T_4334_86;
  wire  T_4334_87;
  wire  T_4334_88;
  wire  T_4334_89;
  wire  T_4334_90;
  wire  T_4334_91;
  wire  T_4334_92;
  wire  T_4334_93;
  wire  T_4334_94;
  wire  T_4334_95;
  wire  T_4334_96;
  wire  T_4334_97;
  wire  T_4334_98;
  wire  T_4334_99;
  wire  T_4334_100;
  wire  T_4334_101;
  wire  T_4334_102;
  wire  T_4334_103;
  wire  T_4334_104;
  wire  T_4334_105;
  wire  T_4334_106;
  wire  T_4334_107;
  wire  T_4334_108;
  wire  T_4334_109;
  wire  T_4334_110;
  wire  T_4334_111;
  wire  T_4334_112;
  wire  T_4334_113;
  wire  T_4334_114;
  wire  T_4334_115;
  wire  T_4334_116;
  wire  T_4334_117;
  wire  T_4334_118;
  wire  T_4334_119;
  wire  T_4334_120;
  wire  T_4334_121;
  wire  T_4334_122;
  wire  T_4334_123;
  wire  T_4334_124;
  wire  T_4334_125;
  wire  T_4334_126;
  wire  T_4334_127;
  wire  T_4334_128;
  wire  T_4334_129;
  wire  T_4334_130;
  wire  T_4334_131;
  wire  T_4334_132;
  wire  T_4334_133;
  wire  T_4334_134;
  wire  T_4334_135;
  wire  T_4334_136;
  wire  T_4334_137;
  wire  T_4334_138;
  wire  T_4334_139;
  wire  T_4334_140;
  wire  T_4334_141;
  wire  T_4334_142;
  wire  T_4334_143;
  wire  T_4334_144;
  wire  T_4334_145;
  wire  T_4334_146;
  wire  T_4334_147;
  wire  T_4334_148;
  wire  T_4334_149;
  wire  T_4334_150;
  wire  T_4334_151;
  wire  T_4334_152;
  wire  T_4334_153;
  wire  T_4334_154;
  wire  T_4334_155;
  wire  T_4334_156;
  wire  T_4334_157;
  wire  T_4339_0;
  wire  T_4339_1;
  wire  T_4339_2;
  wire  T_4339_3;
  wire  T_4339_4;
  wire  T_4339_5;
  wire  T_4339_6;
  wire  T_4339_7;
  wire  T_4339_8;
  wire  T_4339_9;
  wire  T_4339_10;
  wire  T_4339_11;
  wire  T_4339_12;
  wire  T_4339_13;
  wire  T_4339_14;
  wire  T_4339_15;
  wire  T_4339_16;
  wire  T_4339_17;
  wire  T_4339_18;
  wire  T_4339_19;
  wire  T_4339_20;
  wire  T_4339_21;
  wire  T_4339_22;
  wire  T_4339_23;
  wire  T_4339_24;
  wire  T_4339_25;
  wire  T_4339_26;
  wire  T_4339_27;
  wire  T_4339_28;
  wire  T_4339_29;
  wire  T_4339_30;
  wire  T_4339_31;
  wire  T_4339_32;
  wire  T_4339_33;
  wire  T_4339_34;
  wire  T_4339_35;
  wire  T_4339_36;
  wire  T_4339_37;
  wire  T_4339_38;
  wire  T_4339_39;
  wire  T_4339_40;
  wire  T_4339_41;
  wire  T_4339_42;
  wire  T_4339_43;
  wire  T_4339_44;
  wire  T_4339_45;
  wire  T_4339_46;
  wire  T_4339_47;
  wire  T_4339_48;
  wire  T_4339_49;
  wire  T_4339_50;
  wire  T_4339_51;
  wire  T_4339_52;
  wire  T_4339_53;
  wire  T_4339_54;
  wire  T_4339_55;
  wire  T_4339_56;
  wire  T_4339_57;
  wire  T_4339_58;
  wire  T_4339_59;
  wire  T_4339_60;
  wire  T_4339_61;
  wire  T_4339_62;
  wire  T_4339_63;
  wire  T_4339_64;
  wire  T_4339_65;
  wire  T_4339_66;
  wire  T_4339_67;
  wire  T_4339_68;
  wire  T_4339_69;
  wire  T_4339_70;
  wire  T_4339_71;
  wire  T_4339_72;
  wire  T_4339_73;
  wire  T_4339_74;
  wire  T_4339_75;
  wire  T_4339_76;
  wire  T_4339_77;
  wire  T_4339_78;
  wire  T_4339_79;
  wire  T_4339_80;
  wire  T_4339_81;
  wire  T_4339_82;
  wire  T_4339_83;
  wire  T_4339_84;
  wire  T_4339_85;
  wire  T_4339_86;
  wire  T_4339_87;
  wire  T_4339_88;
  wire  T_4339_89;
  wire  T_4339_90;
  wire  T_4339_91;
  wire  T_4339_92;
  wire  T_4339_93;
  wire  T_4339_94;
  wire  T_4339_95;
  wire  T_4339_96;
  wire  T_4339_97;
  wire  T_4339_98;
  wire  T_4339_99;
  wire  T_4339_100;
  wire  T_4339_101;
  wire  T_4339_102;
  wire  T_4339_103;
  wire  T_4339_104;
  wire  T_4339_105;
  wire  T_4339_106;
  wire  T_4339_107;
  wire  T_4339_108;
  wire  T_4339_109;
  wire  T_4339_110;
  wire  T_4339_111;
  wire  T_4339_112;
  wire  T_4339_113;
  wire  T_4339_114;
  wire  T_4339_115;
  wire  T_4339_116;
  wire  T_4339_117;
  wire  T_4339_118;
  wire  T_4339_119;
  wire  T_4339_120;
  wire  T_4339_121;
  wire  T_4339_122;
  wire  T_4339_123;
  wire  T_4339_124;
  wire  T_4339_125;
  wire  T_4339_126;
  wire  T_4339_127;
  wire  T_4339_128;
  wire  T_4339_129;
  wire  T_4339_130;
  wire  T_4339_131;
  wire  T_4339_132;
  wire  T_4339_133;
  wire  T_4339_134;
  wire  T_4339_135;
  wire  T_4339_136;
  wire  T_4339_137;
  wire  T_4339_138;
  wire  T_4339_139;
  wire  T_4339_140;
  wire  T_4339_141;
  wire  T_4339_142;
  wire  T_4339_143;
  wire  T_4339_144;
  wire  T_4339_145;
  wire  T_4339_146;
  wire  T_4339_147;
  wire  T_4339_148;
  wire  T_4339_149;
  wire  T_4339_150;
  wire  T_4339_151;
  wire  T_4339_152;
  wire  T_4339_153;
  wire  T_4339_154;
  wire  T_4339_155;
  wire  T_4339_156;
  wire  T_4339_157;
  wire  T_4344_0;
  wire  T_4344_1;
  wire  T_4344_2;
  wire  T_4344_3;
  wire  T_4344_4;
  wire  T_4344_5;
  wire  T_4344_6;
  wire  T_4344_7;
  wire  T_4344_8;
  wire  T_4344_9;
  wire  T_4344_10;
  wire  T_4344_11;
  wire  T_4344_12;
  wire  T_4344_13;
  wire  T_4344_14;
  wire  T_4344_15;
  wire  T_4344_16;
  wire  T_4344_17;
  wire  T_4344_18;
  wire  T_4344_19;
  wire  T_4344_20;
  wire  T_4344_21;
  wire  T_4344_22;
  wire  T_4344_23;
  wire  T_4344_24;
  wire  T_4344_25;
  wire  T_4344_26;
  wire  T_4344_27;
  wire  T_4344_28;
  wire  T_4344_29;
  wire  T_4344_30;
  wire  T_4344_31;
  wire  T_4344_32;
  wire  T_4344_33;
  wire  T_4344_34;
  wire  T_4344_35;
  wire  T_4344_36;
  wire  T_4344_37;
  wire  T_4344_38;
  wire  T_4344_39;
  wire  T_4344_40;
  wire  T_4344_41;
  wire  T_4344_42;
  wire  T_4344_43;
  wire  T_4344_44;
  wire  T_4344_45;
  wire  T_4344_46;
  wire  T_4344_47;
  wire  T_4344_48;
  wire  T_4344_49;
  wire  T_4344_50;
  wire  T_4344_51;
  wire  T_4344_52;
  wire  T_4344_53;
  wire  T_4344_54;
  wire  T_4344_55;
  wire  T_4344_56;
  wire  T_4344_57;
  wire  T_4344_58;
  wire  T_4344_59;
  wire  T_4344_60;
  wire  T_4344_61;
  wire  T_4344_62;
  wire  T_4344_63;
  wire  T_4344_64;
  wire  T_4344_65;
  wire  T_4344_66;
  wire  T_4344_67;
  wire  T_4344_68;
  wire  T_4344_69;
  wire  T_4344_70;
  wire  T_4344_71;
  wire  T_4344_72;
  wire  T_4344_73;
  wire  T_4344_74;
  wire  T_4344_75;
  wire  T_4344_76;
  wire  T_4344_77;
  wire  T_4344_78;
  wire  T_4344_79;
  wire  T_4344_80;
  wire  T_4344_81;
  wire  T_4344_82;
  wire  T_4344_83;
  wire  T_4344_84;
  wire  T_4344_85;
  wire  T_4344_86;
  wire  T_4344_87;
  wire  T_4344_88;
  wire  T_4344_89;
  wire  T_4344_90;
  wire  T_4344_91;
  wire  T_4344_92;
  wire  T_4344_93;
  wire  T_4344_94;
  wire  T_4344_95;
  wire  T_4344_96;
  wire  T_4344_97;
  wire  T_4344_98;
  wire  T_4344_99;
  wire  T_4344_100;
  wire  T_4344_101;
  wire  T_4344_102;
  wire  T_4344_103;
  wire  T_4344_104;
  wire  T_4344_105;
  wire  T_4344_106;
  wire  T_4344_107;
  wire  T_4344_108;
  wire  T_4344_109;
  wire  T_4344_110;
  wire  T_4344_111;
  wire  T_4344_112;
  wire  T_4344_113;
  wire  T_4344_114;
  wire  T_4344_115;
  wire  T_4344_116;
  wire  T_4344_117;
  wire  T_4344_118;
  wire  T_4344_119;
  wire  T_4344_120;
  wire  T_4344_121;
  wire  T_4344_122;
  wire  T_4344_123;
  wire  T_4344_124;
  wire  T_4344_125;
  wire  T_4344_126;
  wire  T_4344_127;
  wire  T_4344_128;
  wire  T_4344_129;
  wire  T_4344_130;
  wire  T_4344_131;
  wire  T_4344_132;
  wire  T_4344_133;
  wire  T_4344_134;
  wire  T_4344_135;
  wire  T_4344_136;
  wire  T_4344_137;
  wire  T_4344_138;
  wire  T_4344_139;
  wire  T_4344_140;
  wire  T_4344_141;
  wire  T_4344_142;
  wire  T_4344_143;
  wire  T_4344_144;
  wire  T_4344_145;
  wire  T_4344_146;
  wire  T_4344_147;
  wire  T_4344_148;
  wire  T_4344_149;
  wire  T_4344_150;
  wire  T_4344_151;
  wire  T_4344_152;
  wire  T_4344_153;
  wire  T_4344_154;
  wire  T_4344_155;
  wire  T_4344_156;
  wire  T_4344_157;
  wire  T_6906;
  wire  T_6907;
  wire  T_6908;
  wire  T_6909;
  wire [7:0] T_6913;
  wire [7:0] T_6917;
  wire [7:0] T_6921;
  wire [7:0] T_6925;
  wire [15:0] T_6926;
  wire [15:0] T_6927;
  wire [31:0] T_6928;
  wire  T_6952;
  wire  T_6956;
  wire  T_6958;
  wire  T_6972;
  wire  T_6992;
  wire  T_6996;
  wire  T_6998;
  wire  T_7012;
  wire [1:0] GEN_3514;
  wire [1:0] T_7027;
  wire [1:0] GEN_3515;
  wire [1:0] T_7031;
  wire  T_7032;
  wire  T_7036;
  wire  T_7038;
  wire  T_7052;
  wire [2:0] GEN_3516;
  wire [2:0] T_7067;
  wire [2:0] GEN_3517;
  wire [2:0] T_7071;
  wire  T_7072;
  wire  T_7076;
  wire  T_7078;
  wire  T_7092;
  wire [3:0] GEN_3518;
  wire [3:0] T_7107;
  wire [3:0] GEN_3519;
  wire [3:0] T_7111;
  wire  T_7112;
  wire  T_7116;
  wire  T_7118;
  wire  T_7132;
  wire [4:0] GEN_3520;
  wire [4:0] T_7147;
  wire [4:0] GEN_3521;
  wire [4:0] T_7151;
  wire  T_7152;
  wire  T_7156;
  wire  T_7158;
  wire  T_7172;
  wire [5:0] GEN_3522;
  wire [5:0] T_7187;
  wire [5:0] GEN_3523;
  wire [5:0] T_7191;
  wire  T_7192;
  wire  T_7196;
  wire  T_7198;
  wire  T_7212;
  wire [6:0] GEN_3524;
  wire [6:0] T_7227;
  wire [6:0] GEN_3525;
  wire [6:0] T_7231;
  wire  T_7232;
  wire  T_7236;
  wire  T_7238;
  wire  T_7252;
  wire [7:0] GEN_3526;
  wire [7:0] T_7267;
  wire [7:0] GEN_3527;
  wire [7:0] T_7271;
  wire  T_7272;
  wire  T_7276;
  wire  T_7278;
  wire  T_7292;
  wire [8:0] GEN_3528;
  wire [8:0] T_7307;
  wire [8:0] GEN_3529;
  wire [8:0] T_7311;
  wire  T_7312;
  wire  T_7316;
  wire  T_7318;
  wire  T_7332;
  wire [9:0] GEN_3530;
  wire [9:0] T_7347;
  wire [9:0] GEN_3531;
  wire [9:0] T_7351;
  wire  T_7352;
  wire  T_7356;
  wire  T_7358;
  wire  T_7372;
  wire [10:0] GEN_3532;
  wire [10:0] T_7387;
  wire [10:0] GEN_3533;
  wire [10:0] T_7391;
  wire  T_7392;
  wire  T_7396;
  wire  T_7398;
  wire  T_7412;
  wire [11:0] GEN_3534;
  wire [11:0] T_7427;
  wire [11:0] GEN_3535;
  wire [11:0] T_7431;
  wire  T_7432;
  wire  T_7436;
  wire  T_7438;
  wire  T_7452;
  wire [12:0] GEN_3536;
  wire [12:0] T_7467;
  wire [12:0] GEN_3537;
  wire [12:0] T_7471;
  wire  T_7472;
  wire  T_7476;
  wire  T_7478;
  wire  T_7492;
  wire [13:0] GEN_3538;
  wire [13:0] T_7507;
  wire [13:0] GEN_3539;
  wire [13:0] T_7511;
  wire  T_7512;
  wire  T_7516;
  wire  T_7518;
  wire  T_7532;
  wire [14:0] GEN_3540;
  wire [14:0] T_7547;
  wire [14:0] GEN_3541;
  wire [14:0] T_7551;
  wire  T_7552;
  wire  T_7556;
  wire  T_7558;
  wire  T_7572;
  wire [15:0] GEN_3542;
  wire [15:0] T_7587;
  wire [15:0] GEN_3543;
  wire [15:0] T_7591;
  wire  T_7592;
  wire  T_7596;
  wire  T_7598;
  wire  T_7612;
  wire [16:0] GEN_3544;
  wire [16:0] T_7627;
  wire [16:0] GEN_3545;
  wire [16:0] T_7631;
  wire  T_7632;
  wire  T_7636;
  wire  T_7638;
  wire  T_7652;
  wire [17:0] GEN_3546;
  wire [17:0] T_7667;
  wire [17:0] GEN_3547;
  wire [17:0] T_7671;
  wire  T_7672;
  wire  T_7676;
  wire  T_7678;
  wire  T_7692;
  wire [18:0] GEN_3548;
  wire [18:0] T_7707;
  wire [18:0] GEN_3549;
  wire [18:0] T_7711;
  wire  T_7712;
  wire  T_7716;
  wire  T_7718;
  wire  T_7732;
  wire [19:0] GEN_3550;
  wire [19:0] T_7747;
  wire [19:0] GEN_3551;
  wire [19:0] T_7751;
  wire  T_7752;
  wire  T_7756;
  wire  T_7758;
  wire  T_7772;
  wire [20:0] GEN_3552;
  wire [20:0] T_7787;
  wire [20:0] GEN_3553;
  wire [20:0] T_7791;
  wire  T_7792;
  wire  T_7796;
  wire  T_7798;
  wire  T_7812;
  wire [21:0] GEN_3554;
  wire [21:0] T_7827;
  wire [21:0] GEN_3555;
  wire [21:0] T_7831;
  wire  T_7832;
  wire  T_7836;
  wire  T_7838;
  wire  T_7852;
  wire [22:0] GEN_3556;
  wire [22:0] T_7867;
  wire [22:0] GEN_3557;
  wire [22:0] T_7871;
  wire  T_7872;
  wire  T_7876;
  wire  T_7878;
  wire  T_7892;
  wire [23:0] GEN_3558;
  wire [23:0] T_7907;
  wire [23:0] GEN_3559;
  wire [23:0] T_7911;
  wire  T_7912;
  wire  T_7916;
  wire  T_7918;
  wire  T_7932;
  wire [24:0] GEN_3560;
  wire [24:0] T_7947;
  wire [24:0] GEN_3561;
  wire [24:0] T_7951;
  wire  T_7952;
  wire  T_7956;
  wire  T_7958;
  wire  T_7972;
  wire [25:0] GEN_3562;
  wire [25:0] T_7987;
  wire [25:0] GEN_3563;
  wire [25:0] T_7991;
  wire  T_7992;
  wire  T_7996;
  wire  T_7998;
  wire  T_8012;
  wire [26:0] GEN_3564;
  wire [26:0] T_8027;
  wire [26:0] GEN_3565;
  wire [26:0] T_8031;
  wire  T_8032;
  wire  T_8036;
  wire  T_8038;
  wire  T_8052;
  wire [27:0] GEN_3566;
  wire [27:0] T_8067;
  wire [27:0] GEN_3567;
  wire [27:0] T_8071;
  wire  T_8072;
  wire  T_8076;
  wire  T_8078;
  wire  T_8092;
  wire [28:0] GEN_3568;
  wire [28:0] T_8107;
  wire [28:0] GEN_3569;
  wire [28:0] T_8111;
  wire  T_8112;
  wire  T_8116;
  wire  T_8118;
  wire  T_8132;
  wire [29:0] GEN_3570;
  wire [29:0] T_8147;
  wire [29:0] GEN_3571;
  wire [29:0] T_8151;
  wire  T_8152;
  wire  T_8156;
  wire  T_8158;
  wire  T_8172;
  wire [30:0] GEN_3572;
  wire [30:0] T_8187;
  wire [30:0] GEN_3573;
  wire [30:0] T_8191;
  wire  T_8192;
  wire  T_8196;
  wire  T_8198;
  wire  T_8212;
  wire [31:0] GEN_3574;
  wire [31:0] T_8227;
  wire [31:0] GEN_3575;
  wire [31:0] T_8231;
  wire  T_8234;
  wire [31:0] T_8236;
  wire  T_8238;
  wire [31:0] T_8270;
  wire  T_8291;
  wire [31:0] GEN_61;
  wire [31:0] T_8310;
  wire  T_8331;
  wire [31:0] GEN_62;
  wire [31:0] T_8350;
  wire  T_8371;
  wire [31:0] GEN_63;
  wire [31:0] T_8390;
  wire  T_8411;
  wire [31:0] GEN_64;
  wire [31:0] T_8430;
  wire  T_8451;
  wire [31:0] GEN_65;
  wire [31:0] T_8470;
  wire  T_8491;
  wire [31:0] GEN_66;
  wire [31:0] T_8510;
  wire  T_8531;
  wire [31:0] GEN_67;
  wire [31:0] T_8550;
  wire  T_8571;
  wire [31:0] GEN_68;
  wire [31:0] T_8590;
  wire  T_8611;
  wire  GEN_69;
  wire  T_8651;
  wire  GEN_70;
  wire [1:0] GEN_3576;
  wire [1:0] T_8667;
  wire [1:0] GEN_3577;
  wire [1:0] T_8671;
  wire  T_8691;
  wire  GEN_71;
  wire [2:0] GEN_3578;
  wire [2:0] T_8707;
  wire [2:0] GEN_3579;
  wire [2:0] T_8711;
  wire  T_8731;
  wire  GEN_72;
  wire [3:0] GEN_3580;
  wire [3:0] T_8747;
  wire [3:0] GEN_3581;
  wire [3:0] T_8751;
  wire  T_8771;
  wire  GEN_73;
  wire [4:0] GEN_3582;
  wire [4:0] T_8787;
  wire [4:0] GEN_3583;
  wire [4:0] T_8791;
  wire  T_8811;
  wire  GEN_74;
  wire [5:0] GEN_3584;
  wire [5:0] T_8827;
  wire [5:0] GEN_3585;
  wire [5:0] T_8831;
  wire  T_8851;
  wire  GEN_75;
  wire [6:0] GEN_3586;
  wire [6:0] T_8867;
  wire [6:0] GEN_3587;
  wire [6:0] T_8871;
  wire  T_8891;
  wire  GEN_76;
  wire [7:0] GEN_3588;
  wire [7:0] T_8907;
  wire [7:0] GEN_3589;
  wire [7:0] T_8911;
  wire  T_8931;
  wire  GEN_77;
  wire [8:0] GEN_3590;
  wire [8:0] T_8947;
  wire [8:0] GEN_3591;
  wire [8:0] T_8951;
  wire  T_8971;
  wire  GEN_78;
  wire [9:0] GEN_3592;
  wire [9:0] T_8987;
  wire [9:0] GEN_3593;
  wire [9:0] T_8991;
  wire  T_9011;
  wire  GEN_79;
  wire [10:0] GEN_3594;
  wire [10:0] T_9027;
  wire [10:0] GEN_3595;
  wire [10:0] T_9031;
  wire  T_9051;
  wire  GEN_80;
  wire [11:0] GEN_3596;
  wire [11:0] T_9067;
  wire [11:0] GEN_3597;
  wire [11:0] T_9071;
  wire  T_9091;
  wire  GEN_81;
  wire [12:0] GEN_3598;
  wire [12:0] T_9107;
  wire [12:0] GEN_3599;
  wire [12:0] T_9111;
  wire  T_9131;
  wire  GEN_82;
  wire [13:0] GEN_3600;
  wire [13:0] T_9147;
  wire [13:0] GEN_3601;
  wire [13:0] T_9151;
  wire  T_9171;
  wire  GEN_83;
  wire [14:0] GEN_3602;
  wire [14:0] T_9187;
  wire [14:0] GEN_3603;
  wire [14:0] T_9191;
  wire  T_9211;
  wire  GEN_84;
  wire [15:0] GEN_3604;
  wire [15:0] T_9227;
  wire [15:0] GEN_3605;
  wire [15:0] T_9231;
  wire  T_9251;
  wire  GEN_85;
  wire [16:0] GEN_3606;
  wire [16:0] T_9267;
  wire [16:0] GEN_3607;
  wire [16:0] T_9271;
  wire  T_9291;
  wire  GEN_86;
  wire [17:0] GEN_3608;
  wire [17:0] T_9307;
  wire [17:0] GEN_3609;
  wire [17:0] T_9311;
  wire  T_9331;
  wire  GEN_87;
  wire [18:0] GEN_3610;
  wire [18:0] T_9347;
  wire [18:0] GEN_3611;
  wire [18:0] T_9351;
  wire  T_9371;
  wire  GEN_88;
  wire [19:0] GEN_3612;
  wire [19:0] T_9387;
  wire [19:0] GEN_3613;
  wire [19:0] T_9391;
  wire  T_9411;
  wire [31:0] GEN_89;
  wire [31:0] T_9430;
  wire  T_9451;
  wire [31:0] GEN_90;
  wire [31:0] T_9470;
  wire  T_9487;
  wire  GEN_0;
  wire  GEN_92;
  wire  GEN_93;
  wire  GEN_94;
  wire  GEN_95;
  wire  GEN_96;
  wire  GEN_97;
  wire  GEN_98;
  wire  GEN_99;
  wire  GEN_100;
  wire  GEN_101;
  wire  GEN_102;
  wire  GEN_103;
  wire  GEN_104;
  wire  GEN_105;
  wire  GEN_106;
  wire  GEN_107;
  wire  GEN_108;
  wire  GEN_109;
  wire  GEN_110;
  wire  GEN_111;
  wire  GEN_112;
  wire  GEN_113;
  wire  GEN_114;
  wire  GEN_115;
  wire  GEN_116;
  wire  GEN_117;
  wire  GEN_118;
  wire  GEN_119;
  wire  GEN_120;
  wire  GEN_121;
  wire  GEN_122;
  wire  GEN_123;
  wire  GEN_124;
  wire  GEN_125;
  wire  GEN_126;
  wire  GEN_127;
  wire  GEN_128;
  wire  GEN_129;
  wire  GEN_130;
  wire  GEN_131;
  wire  GEN_132;
  wire  GEN_133;
  wire  GEN_134;
  wire  GEN_135;
  wire  GEN_136;
  wire  GEN_137;
  wire  GEN_138;
  wire  GEN_139;
  wire  GEN_140;
  wire  GEN_141;
  wire  GEN_142;
  wire  GEN_144;
  wire  GEN_145;
  wire  GEN_146;
  wire  GEN_147;
  wire  GEN_148;
  wire  GEN_149;
  wire  GEN_150;
  wire  GEN_151;
  wire  GEN_152;
  wire  GEN_153;
  wire  GEN_154;
  wire  GEN_155;
  wire  GEN_156;
  wire  GEN_157;
  wire  GEN_158;
  wire  GEN_159;
  wire  GEN_160;
  wire  GEN_161;
  wire  GEN_162;
  wire  GEN_163;
  wire  GEN_164;
  wire  GEN_165;
  wire  GEN_166;
  wire  GEN_167;
  wire  GEN_168;
  wire  GEN_169;
  wire  GEN_170;
  wire  GEN_171;
  wire  GEN_172;
  wire  GEN_173;
  wire  GEN_174;
  wire  GEN_175;
  wire  GEN_176;
  wire  GEN_177;
  wire  GEN_178;
  wire  GEN_179;
  wire  GEN_180;
  wire  GEN_181;
  wire  GEN_182;
  wire  GEN_183;
  wire  GEN_184;
  wire  GEN_185;
  wire  GEN_186;
  wire  GEN_187;
  wire  GEN_188;
  wire  GEN_189;
  wire  GEN_190;
  wire  GEN_191;
  wire  GEN_192;
  wire  GEN_193;
  wire  GEN_194;
  wire [5:0] GEN_195;
  wire  T_9494;
  wire [5:0] T_9497;
  wire  GEN_1;
  wire  GEN_196;
  wire  GEN_197;
  wire  GEN_198;
  wire  GEN_199;
  wire  GEN_200;
  wire  GEN_201;
  wire  GEN_202;
  wire  GEN_203;
  wire  GEN_204;
  wire  GEN_205;
  wire  GEN_206;
  wire  GEN_207;
  wire  GEN_208;
  wire  GEN_209;
  wire  GEN_210;
  wire  GEN_211;
  wire  GEN_212;
  wire  GEN_213;
  wire  GEN_214;
  wire  GEN_215;
  wire  GEN_216;
  wire  GEN_217;
  wire  GEN_218;
  wire  GEN_219;
  wire  GEN_220;
  wire  GEN_221;
  wire  GEN_222;
  wire  GEN_223;
  wire  GEN_224;
  wire  GEN_225;
  wire  GEN_226;
  wire  GEN_227;
  wire  GEN_228;
  wire  GEN_229;
  wire  GEN_230;
  wire  GEN_231;
  wire  GEN_232;
  wire  GEN_233;
  wire  GEN_234;
  wire  GEN_235;
  wire  GEN_236;
  wire  GEN_237;
  wire  GEN_238;
  wire  GEN_239;
  wire  GEN_240;
  wire  GEN_241;
  wire  GEN_242;
  wire  GEN_243;
  wire  GEN_244;
  wire  GEN_245;
  wire  GEN_246;
  wire  T_9498;
  wire [32:0] T_9500;
  wire [31:0] T_9501;
  wire [5:0] T_9515;
  wire  GEN_2;
  wire  GEN_247;
  wire  GEN_248;
  wire  GEN_249;
  wire  GEN_250;
  wire  GEN_251;
  wire  GEN_252;
  wire  GEN_253;
  wire  GEN_254;
  wire  GEN_255;
  wire  GEN_256;
  wire  GEN_257;
  wire  GEN_258;
  wire  GEN_259;
  wire  GEN_260;
  wire  GEN_261;
  wire  GEN_262;
  wire  GEN_263;
  wire  GEN_264;
  wire  GEN_265;
  wire  GEN_266;
  wire  GEN_267;
  wire  GEN_268;
  wire  GEN_269;
  wire  GEN_270;
  wire  GEN_271;
  wire  GEN_272;
  wire  GEN_273;
  wire  GEN_274;
  wire  GEN_275;
  wire  GEN_276;
  wire  GEN_277;
  wire  GEN_278;
  wire  GEN_279;
  wire  GEN_280;
  wire  GEN_281;
  wire  GEN_282;
  wire  GEN_283;
  wire  GEN_284;
  wire  GEN_285;
  wire  GEN_286;
  wire  GEN_287;
  wire  GEN_288;
  wire  GEN_289;
  wire  GEN_290;
  wire  GEN_291;
  wire  GEN_292;
  wire  GEN_293;
  wire  GEN_294;
  wire  GEN_295;
  wire  GEN_296;
  wire  GEN_297;
  wire  GEN_298;
  wire  GEN_299;
  wire  GEN_300;
  wire  GEN_301;
  wire  GEN_302;
  wire  GEN_303;
  wire  GEN_304;
  wire  GEN_305;
  wire  GEN_306;
  wire  GEN_307;
  wire  GEN_308;
  wire  GEN_309;
  wire  GEN_310;
  wire  GEN_311;
  wire  GEN_312;
  wire  GEN_313;
  wire  GEN_314;
  wire  GEN_315;
  wire  GEN_316;
  wire  GEN_317;
  wire  GEN_318;
  wire  GEN_319;
  wire  GEN_320;
  wire  GEN_321;
  wire  GEN_322;
  wire  GEN_323;
  wire  GEN_324;
  wire  GEN_325;
  wire  GEN_326;
  wire  GEN_327;
  wire  GEN_328;
  wire  GEN_329;
  wire  GEN_330;
  wire  GEN_331;
  wire  GEN_332;
  wire  GEN_333;
  wire  GEN_334;
  wire  GEN_335;
  wire  GEN_336;
  wire  GEN_337;
  wire  GEN_338;
  wire  GEN_339;
  wire  GEN_340;
  wire  GEN_341;
  wire  GEN_342;
  wire  GEN_343;
  wire  GEN_344;
  wire  GEN_345;
  wire  GEN_346;
  wire  GEN_347;
  wire  GEN_348;
  wire [31:0] T_9533;
  wire  T_9554;
  wire [31:0] GEN_349;
  wire [31:0] T_9573;
  wire  T_9594;
  wire [31:0] GEN_350;
  wire [31:0] T_9613;
  wire  T_9634;
  wire [31:0] GEN_351;
  wire [31:0] T_9653;
  wire  T_9674;
  wire [31:0] GEN_352;
  wire [31:0] T_9693;
  wire  T_9714;
  wire [31:0] GEN_353;
  wire [31:0] T_9733;
  wire  T_9754;
  wire [31:0] GEN_354;
  wire [31:0] T_9773;
  wire  T_9794;
  wire [31:0] GEN_355;
  wire [31:0] T_9813;
  wire  T_9834;
  wire [31:0] GEN_356;
  wire [31:0] T_9853;
  wire  T_9874;
  wire [31:0] GEN_357;
  wire [31:0] T_9893;
  wire  T_9914;
  wire [31:0] GEN_358;
  wire [31:0] T_9933;
  wire  T_9954;
  wire [31:0] GEN_359;
  wire [31:0] T_9973;
  wire  T_9994;
  wire [31:0] GEN_360;
  wire [31:0] T_10013;
  wire  T_10034;
  wire [31:0] GEN_361;
  wire [31:0] T_10053;
  wire  T_10074;
  wire [31:0] GEN_362;
  wire [31:0] T_10093;
  wire  T_10114;
  wire [31:0] GEN_363;
  wire [31:0] T_10133;
  wire  T_10194;
  wire  GEN_365;
  wire [1:0] GEN_3614;
  wire [1:0] T_10210;
  wire [1:0] GEN_3615;
  wire [1:0] T_10214;
  wire  T_10234;
  wire  GEN_366;
  wire [2:0] GEN_3616;
  wire [2:0] T_10250;
  wire [2:0] GEN_3617;
  wire [2:0] T_10254;
  wire  T_10274;
  wire  GEN_367;
  wire [3:0] GEN_3618;
  wire [3:0] T_10290;
  wire [3:0] GEN_3619;
  wire [3:0] T_10294;
  wire  T_10314;
  wire  GEN_368;
  wire [4:0] GEN_3620;
  wire [4:0] T_10330;
  wire [4:0] GEN_3621;
  wire [4:0] T_10334;
  wire  T_10354;
  wire  GEN_369;
  wire [5:0] GEN_3622;
  wire [5:0] T_10370;
  wire [5:0] GEN_3623;
  wire [5:0] T_10374;
  wire  T_10394;
  wire  GEN_370;
  wire [6:0] GEN_3624;
  wire [6:0] T_10410;
  wire [6:0] GEN_3625;
  wire [6:0] T_10414;
  wire  T_10434;
  wire  GEN_371;
  wire [7:0] GEN_3626;
  wire [7:0] T_10450;
  wire [7:0] GEN_3627;
  wire [7:0] T_10454;
  wire  T_10474;
  wire  GEN_372;
  wire [8:0] GEN_3628;
  wire [8:0] T_10490;
  wire [8:0] GEN_3629;
  wire [8:0] T_10494;
  wire  T_10514;
  wire  GEN_373;
  wire [9:0] GEN_3630;
  wire [9:0] T_10530;
  wire [9:0] GEN_3631;
  wire [9:0] T_10534;
  wire  T_10554;
  wire  GEN_374;
  wire [10:0] GEN_3632;
  wire [10:0] T_10570;
  wire [10:0] GEN_3633;
  wire [10:0] T_10574;
  wire  T_10594;
  wire  GEN_375;
  wire [11:0] GEN_3634;
  wire [11:0] T_10610;
  wire [11:0] GEN_3635;
  wire [11:0] T_10614;
  wire  T_10634;
  wire  GEN_376;
  wire [12:0] GEN_3636;
  wire [12:0] T_10650;
  wire [12:0] GEN_3637;
  wire [12:0] T_10654;
  wire  T_10674;
  wire  GEN_377;
  wire [13:0] GEN_3638;
  wire [13:0] T_10690;
  wire [13:0] GEN_3639;
  wire [13:0] T_10694;
  wire  T_10714;
  wire  GEN_378;
  wire [14:0] GEN_3640;
  wire [14:0] T_10730;
  wire [14:0] GEN_3641;
  wire [14:0] T_10734;
  wire  T_10754;
  wire  GEN_379;
  wire [15:0] GEN_3642;
  wire [15:0] T_10770;
  wire [15:0] GEN_3643;
  wire [15:0] T_10774;
  wire  T_10794;
  wire  GEN_380;
  wire [16:0] GEN_3644;
  wire [16:0] T_10810;
  wire [16:0] GEN_3645;
  wire [16:0] T_10814;
  wire  T_10834;
  wire  GEN_381;
  wire [17:0] GEN_3646;
  wire [17:0] T_10850;
  wire [17:0] GEN_3647;
  wire [17:0] T_10854;
  wire  T_10874;
  wire  GEN_382;
  wire [18:0] GEN_3648;
  wire [18:0] T_10890;
  wire [18:0] GEN_3649;
  wire [18:0] T_10894;
  wire  T_10914;
  wire  GEN_383;
  wire [19:0] GEN_3650;
  wire [19:0] T_10930;
  wire [19:0] GEN_3651;
  wire [19:0] T_10934;
  wire  T_10954;
  wire  GEN_384;
  wire [20:0] GEN_3652;
  wire [20:0] T_10970;
  wire [20:0] GEN_3653;
  wire [20:0] T_10974;
  wire  T_10994;
  wire  GEN_385;
  wire [21:0] GEN_3654;
  wire [21:0] T_11010;
  wire [21:0] GEN_3655;
  wire [21:0] T_11014;
  wire  T_11034;
  wire  GEN_386;
  wire [22:0] GEN_3656;
  wire [22:0] T_11050;
  wire [22:0] GEN_3657;
  wire [22:0] T_11054;
  wire  T_11074;
  wire  GEN_387;
  wire [23:0] GEN_3658;
  wire [23:0] T_11090;
  wire [23:0] GEN_3659;
  wire [23:0] T_11094;
  wire  T_11114;
  wire  GEN_388;
  wire [24:0] GEN_3660;
  wire [24:0] T_11130;
  wire [24:0] GEN_3661;
  wire [24:0] T_11134;
  wire  T_11154;
  wire  GEN_389;
  wire [25:0] GEN_3662;
  wire [25:0] T_11170;
  wire [25:0] GEN_3663;
  wire [25:0] T_11174;
  wire  T_11194;
  wire  GEN_390;
  wire [26:0] GEN_3664;
  wire [26:0] T_11210;
  wire [26:0] GEN_3665;
  wire [26:0] T_11214;
  wire  T_11234;
  wire  GEN_391;
  wire [27:0] GEN_3666;
  wire [27:0] T_11250;
  wire [27:0] GEN_3667;
  wire [27:0] T_11254;
  wire  T_11274;
  wire  GEN_392;
  wire [28:0] GEN_3668;
  wire [28:0] T_11290;
  wire [28:0] GEN_3669;
  wire [28:0] T_11294;
  wire  T_11314;
  wire  GEN_393;
  wire [29:0] GEN_3670;
  wire [29:0] T_11330;
  wire [29:0] GEN_3671;
  wire [29:0] T_11334;
  wire  T_11354;
  wire  GEN_394;
  wire [30:0] GEN_3672;
  wire [30:0] T_11370;
  wire [30:0] GEN_3673;
  wire [30:0] T_11374;
  wire  T_11394;
  wire  GEN_395;
  wire [31:0] GEN_3674;
  wire [31:0] T_11410;
  wire [31:0] GEN_3675;
  wire [31:0] T_11414;
  wire  T_11434;
  wire [31:0] GEN_396;
  wire [31:0] T_11453;
  wire  T_11474;
  wire [31:0] GEN_397;
  wire [31:0] T_11493;
  wire  T_11514;
  wire [31:0] GEN_398;
  wire [31:0] T_11533;
  wire  T_11554;
  wire [31:0] GEN_399;
  wire [31:0] T_11573;
  wire  T_11594;
  wire [31:0] GEN_400;
  wire [31:0] T_11613;
  wire  T_11634;
  wire [31:0] GEN_401;
  wire [31:0] T_11653;
  wire  T_11674;
  wire [31:0] GEN_402;
  wire [31:0] T_11693;
  wire  T_11714;
  wire [31:0] GEN_403;
  wire [31:0] T_11733;
  wire  T_11754;
  wire [31:0] GEN_404;
  wire [31:0] T_11773;
  wire  T_11794;
  wire [31:0] GEN_405;
  wire [31:0] T_11813;
  wire [1:0] GEN_3676;
  wire [1:0] T_11890;
  wire [1:0] GEN_3677;
  wire [1:0] T_11894;
  wire [2:0] GEN_3678;
  wire [2:0] T_11930;
  wire [2:0] GEN_3679;
  wire [2:0] T_11934;
  wire [3:0] GEN_3680;
  wire [3:0] T_11970;
  wire [3:0] GEN_3681;
  wire [3:0] T_11974;
  wire [4:0] GEN_3682;
  wire [4:0] T_12010;
  wire [4:0] GEN_3683;
  wire [4:0] T_12014;
  wire [5:0] GEN_3684;
  wire [5:0] T_12050;
  wire [5:0] GEN_3685;
  wire [5:0] T_12054;
  wire [6:0] GEN_3686;
  wire [6:0] T_12090;
  wire [6:0] GEN_3687;
  wire [6:0] T_12094;
  wire [7:0] GEN_3688;
  wire [7:0] T_12130;
  wire [7:0] GEN_3689;
  wire [7:0] T_12134;
  wire [8:0] GEN_3690;
  wire [8:0] T_12170;
  wire [8:0] GEN_3691;
  wire [8:0] T_12174;
  wire [9:0] GEN_3692;
  wire [9:0] T_12210;
  wire [9:0] GEN_3693;
  wire [9:0] T_12214;
  wire [10:0] GEN_3694;
  wire [10:0] T_12250;
  wire [10:0] GEN_3695;
  wire [10:0] T_12254;
  wire [11:0] GEN_3696;
  wire [11:0] T_12290;
  wire [11:0] GEN_3697;
  wire [11:0] T_12294;
  wire [12:0] GEN_3698;
  wire [12:0] T_12330;
  wire [12:0] GEN_3699;
  wire [12:0] T_12334;
  wire [13:0] GEN_3700;
  wire [13:0] T_12370;
  wire [13:0] GEN_3701;
  wire [13:0] T_12374;
  wire [14:0] GEN_3702;
  wire [14:0] T_12410;
  wire [14:0] GEN_3703;
  wire [14:0] T_12414;
  wire [15:0] GEN_3704;
  wire [15:0] T_12450;
  wire [15:0] GEN_3705;
  wire [15:0] T_12454;
  wire [16:0] GEN_3706;
  wire [16:0] T_12490;
  wire [16:0] GEN_3707;
  wire [16:0] T_12494;
  wire [17:0] GEN_3708;
  wire [17:0] T_12530;
  wire [17:0] GEN_3709;
  wire [17:0] T_12534;
  wire [18:0] GEN_3710;
  wire [18:0] T_12570;
  wire [18:0] GEN_3711;
  wire [18:0] T_12574;
  wire [19:0] GEN_3712;
  wire [19:0] T_12610;
  wire [19:0] GEN_3713;
  wire [19:0] T_12614;
  wire  T_12634;
  wire [31:0] GEN_406;
  wire [31:0] T_12653;
  wire  T_12674;
  wire [31:0] GEN_407;
  wire [31:0] T_12693;
  wire  T_12714;
  wire [31:0] GEN_408;
  wire [31:0] T_12733;
  wire  T_12754;
  wire [31:0] GEN_409;
  wire [31:0] T_12773;
  wire  T_12794;
  wire [31:0] GEN_410;
  wire [31:0] T_12813;
  wire  T_12834;
  wire [31:0] GEN_411;
  wire [31:0] T_12853;
  wire  T_12874;
  wire [31:0] GEN_412;
  wire [31:0] T_12893;
  wire  T_12914;
  wire [31:0] GEN_413;
  wire [31:0] T_12933;
  wire  T_12954;
  wire [31:0] GEN_414;
  wire [31:0] T_12973;
  wire  T_12994;
  wire [31:0] GEN_415;
  wire [31:0] T_13013;
  wire  T_13034;
  wire [31:0] GEN_416;
  wire [31:0] T_13053;
  wire  T_13074;
  wire [31:0] GEN_417;
  wire [31:0] T_13093;
  wire  T_13114;
  wire [31:0] GEN_418;
  wire [31:0] T_13133;
  wire  T_13154;
  wire [31:0] GEN_419;
  wire [31:0] T_13173;
  wire  T_13194;
  wire [31:0] GEN_420;
  wire [31:0] T_13213;
  wire  T_13234;
  wire [31:0] GEN_421;
  wire [31:0] T_13253;
  wire  T_13274;
  wire [31:0] GEN_422;
  wire [31:0] T_13293;
  wire  T_13541;
  wire  T_13542;
  wire  T_13543;
  wire  T_13544;
  wire  T_13545;
  wire  T_13546;
  wire  T_13547;
  wire  T_13548;
  wire  T_13549;
  wire  T_13550;
  wire  T_13551;
  wire  T_13552;
  wire  T_13553;
  wire  T_13554;
  wire  T_13555;
  wire  T_13556;
  wire  T_13557;
  wire  T_13558;
  wire  T_13559;
  wire  T_13560;
  wire  T_13561;
  wire  T_13562;
  wire  T_13563;
  wire  T_13564;
  wire  T_13565;
  wire  T_13566;
  wire  T_13567;
  wire  T_13568;
  wire  T_13569;
  wire  T_13570;
  wire  T_13571;
  wire  T_13576;
  wire  T_13577;
  wire  T_13578;
  wire  T_13579;
  wire  T_13580;
  wire  T_13581;
  wire  T_13582;
  wire  T_13583;
  wire  T_13584;
  wire  T_13585;
  wire  T_13586;
  wire  T_13587;
  wire  T_13588;
  wire  T_13589;
  wire  T_13590;
  wire  T_13591;
  wire  T_13592;
  wire  T_13593;
  wire  T_13594;
  wire  T_13785;
  wire  T_13786;
  wire  T_13787;
  wire  T_13788;
  wire  T_13789;
  wire  T_13790;
  wire  T_13791;
  wire  T_13792;
  wire  T_13793;
  wire  T_13794;
  wire  T_13795;
  wire  T_13796;
  wire  T_13797;
  wire  T_13798;
  wire  T_13799;
  wire  T_13800;
  wire  T_13801;
  wire  T_13802;
  wire  T_13803;
  wire  T_13804;
  wire  T_13805;
  wire  T_13806;
  wire  T_13807;
  wire  T_13808;
  wire  T_13809;
  wire  T_13810;
  wire  T_13811;
  wire  T_13812;
  wire  T_13813;
  wire  T_13814;
  wire  T_13815;
  wire  T_13820;
  wire  T_13821;
  wire  T_13822;
  wire  T_13823;
  wire  T_13824;
  wire  T_13825;
  wire  T_13826;
  wire  T_13827;
  wire  T_13828;
  wire  T_13829;
  wire  T_13830;
  wire  T_13831;
  wire  T_13832;
  wire  T_13833;
  wire  T_13834;
  wire  T_13835;
  wire  T_13836;
  wire  T_13837;
  wire  T_13838;
  wire  T_15504_0;
  wire  T_15504_1;
  wire  T_15504_2;
  wire  T_15504_3;
  wire  T_15504_4;
  wire  T_15504_5;
  wire  T_15504_6;
  wire  T_15504_7;
  wire  T_15504_8;
  wire  T_15504_9;
  wire  T_15504_10;
  wire  T_15504_11;
  wire  T_15504_12;
  wire  T_15504_13;
  wire  T_15504_14;
  wire  T_15504_15;
  wire  T_15504_16;
  wire  T_15504_17;
  wire  T_15504_18;
  wire  T_15504_19;
  wire  T_15504_20;
  wire  T_15504_21;
  wire  T_15504_22;
  wire  T_15504_23;
  wire  T_15504_24;
  wire  T_15504_25;
  wire  T_15504_26;
  wire  T_15504_27;
  wire  T_15504_28;
  wire  T_15504_29;
  wire  T_15504_30;
  wire  T_15504_31;
  wire  T_15504_32;
  wire  T_15504_33;
  wire  T_15504_34;
  wire  T_15504_35;
  wire  T_15504_36;
  wire  T_15504_37;
  wire  T_15504_38;
  wire  T_15504_39;
  wire  T_15504_40;
  wire  T_15504_41;
  wire  T_15504_42;
  wire  T_15504_43;
  wire  T_15504_44;
  wire  T_15504_45;
  wire  T_15504_46;
  wire  T_15504_47;
  wire  T_15504_48;
  wire  T_15504_49;
  wire  T_15504_50;
  wire  T_15504_51;
  wire  T_15504_52;
  wire  T_15504_53;
  wire  T_15504_54;
  wire  T_15504_55;
  wire  T_15504_56;
  wire  T_15504_57;
  wire  T_15504_58;
  wire  T_15504_59;
  wire  T_15504_60;
  wire  T_15504_61;
  wire  T_15504_62;
  wire  T_15504_63;
  wire  T_15504_64;
  wire  T_15504_65;
  wire  T_15504_66;
  wire  T_15504_67;
  wire  T_15504_68;
  wire  T_15504_69;
  wire  T_15504_70;
  wire  T_15504_71;
  wire  T_15504_72;
  wire  T_15504_73;
  wire  T_15504_74;
  wire  T_15504_75;
  wire  T_15504_76;
  wire  T_15504_77;
  wire  T_15504_78;
  wire  T_15504_79;
  wire  T_15504_80;
  wire  T_15504_81;
  wire  T_15504_82;
  wire  T_15504_83;
  wire  T_15504_84;
  wire  T_15504_85;
  wire  T_15504_86;
  wire  T_15504_87;
  wire  T_15504_88;
  wire  T_15504_89;
  wire  T_15504_90;
  wire  T_15504_91;
  wire  T_15504_92;
  wire  T_15504_93;
  wire  T_15504_94;
  wire  T_15504_95;
  wire  T_15504_96;
  wire  T_15504_97;
  wire  T_15504_98;
  wire  T_15504_99;
  wire  T_15504_100;
  wire  T_15504_101;
  wire  T_15504_102;
  wire  T_15504_103;
  wire  T_15504_104;
  wire  T_15504_105;
  wire  T_15504_106;
  wire  T_15504_107;
  wire  T_15504_108;
  wire  T_15504_109;
  wire  T_15504_110;
  wire  T_15504_111;
  wire  T_15504_112;
  wire  T_15504_113;
  wire  T_15504_114;
  wire  T_15504_115;
  wire  T_15504_116;
  wire  T_15504_117;
  wire  T_15504_118;
  wire  T_15504_119;
  wire  T_15504_120;
  wire  T_15504_121;
  wire  T_15504_122;
  wire  T_15504_123;
  wire  T_15504_124;
  wire  T_15504_125;
  wire  T_15504_126;
  wire  T_15504_127;
  wire  T_15504_128;
  wire  T_15504_129;
  wire  T_15504_130;
  wire  T_15504_131;
  wire  T_15504_132;
  wire  T_15504_133;
  wire  T_15504_134;
  wire  T_15504_135;
  wire  T_15504_136;
  wire  T_15504_137;
  wire  T_15504_138;
  wire  T_15504_139;
  wire  T_15504_140;
  wire  T_15504_141;
  wire  T_15504_142;
  wire  T_15504_143;
  wire  T_15504_144;
  wire  T_15504_145;
  wire  T_15504_146;
  wire  T_15504_147;
  wire  T_15504_148;
  wire  T_15504_149;
  wire  T_15504_150;
  wire  T_15504_151;
  wire  T_15504_152;
  wire  T_15504_153;
  wire  T_15504_154;
  wire  T_15504_155;
  wire  T_15504_156;
  wire  T_15504_157;
  wire  T_15504_158;
  wire  T_15504_159;
  wire  T_15504_160;
  wire  T_15504_161;
  wire  T_15504_162;
  wire  T_15504_163;
  wire  T_15504_164;
  wire  T_15504_165;
  wire  T_15504_166;
  wire  T_15504_167;
  wire  T_15504_168;
  wire  T_15504_169;
  wire  T_15504_170;
  wire  T_15504_171;
  wire  T_15504_172;
  wire  T_15504_173;
  wire  T_15504_174;
  wire  T_15504_175;
  wire  T_15504_176;
  wire  T_15504_177;
  wire  T_15504_178;
  wire  T_15504_179;
  wire  T_15504_180;
  wire  T_15504_181;
  wire  T_15504_182;
  wire  T_15504_183;
  wire  T_15504_184;
  wire  T_15504_185;
  wire  T_15504_186;
  wire  T_15504_187;
  wire  T_15504_188;
  wire  T_15504_189;
  wire  T_15504_190;
  wire  T_15504_191;
  wire  T_15504_192;
  wire  T_15504_193;
  wire  T_15504_194;
  wire  T_15504_195;
  wire  T_15504_196;
  wire  T_15504_197;
  wire  T_15504_198;
  wire  T_15504_199;
  wire  T_15504_200;
  wire  T_15504_201;
  wire  T_15504_202;
  wire  T_15504_203;
  wire  T_15504_204;
  wire  T_15504_205;
  wire  T_15504_206;
  wire  T_15504_207;
  wire  T_15504_208;
  wire  T_15504_209;
  wire  T_15504_210;
  wire  T_15504_211;
  wire  T_15504_212;
  wire  T_15504_213;
  wire  T_15504_214;
  wire  T_15504_215;
  wire  T_15504_216;
  wire  T_15504_217;
  wire  T_15504_218;
  wire  T_15504_219;
  wire  T_15504_220;
  wire  T_15504_221;
  wire  T_15504_222;
  wire  T_15504_223;
  wire  T_15504_224;
  wire  T_15504_225;
  wire  T_15504_226;
  wire  T_15504_227;
  wire  T_15504_228;
  wire  T_15504_229;
  wire  T_15504_230;
  wire  T_15504_231;
  wire  T_15504_232;
  wire  T_15504_233;
  wire  T_15504_234;
  wire  T_15504_235;
  wire  T_15504_236;
  wire  T_15504_237;
  wire  T_15504_238;
  wire  T_15504_239;
  wire  T_15504_240;
  wire  T_15504_241;
  wire  T_15504_242;
  wire  T_15504_243;
  wire  T_15504_244;
  wire  T_15504_245;
  wire  T_15504_246;
  wire  T_15504_247;
  wire  T_15504_248;
  wire  T_15504_249;
  wire  T_15504_250;
  wire  T_15504_251;
  wire  T_15504_252;
  wire  T_15504_253;
  wire  T_15504_254;
  wire  T_15504_255;
  wire  T_15504_256;
  wire  T_15504_257;
  wire  T_15504_258;
  wire  T_15504_259;
  wire  T_15504_260;
  wire  T_15504_261;
  wire  T_15504_262;
  wire  T_15504_263;
  wire  T_15504_264;
  wire  T_15504_265;
  wire  T_15504_266;
  wire  T_15504_267;
  wire  T_15504_268;
  wire  T_15504_269;
  wire  T_15504_270;
  wire  T_15504_271;
  wire  T_15504_272;
  wire  T_15504_273;
  wire  T_15504_274;
  wire  T_15504_275;
  wire  T_15504_276;
  wire  T_15504_277;
  wire  T_15504_278;
  wire  T_15504_279;
  wire  T_15504_280;
  wire  T_15504_281;
  wire  T_15504_282;
  wire  T_15504_283;
  wire  T_15504_284;
  wire  T_15504_285;
  wire  T_15504_286;
  wire  T_15504_287;
  wire  T_15504_288;
  wire  T_15504_289;
  wire  T_15504_290;
  wire  T_15504_291;
  wire  T_15504_292;
  wire  T_15504_293;
  wire  T_15504_294;
  wire  T_15504_295;
  wire  T_15504_296;
  wire  T_15504_297;
  wire  T_15504_298;
  wire  T_15504_299;
  wire  T_15504_300;
  wire  T_15504_301;
  wire  T_15504_302;
  wire  T_15504_303;
  wire  T_15504_304;
  wire  T_15504_305;
  wire  T_15504_306;
  wire  T_15504_307;
  wire  T_15504_308;
  wire  T_15504_309;
  wire  T_15504_310;
  wire  T_15504_311;
  wire  T_15504_312;
  wire  T_15504_313;
  wire  T_15504_314;
  wire  T_15504_315;
  wire  T_15504_316;
  wire  T_15504_317;
  wire  T_15504_318;
  wire  T_15504_319;
  wire  T_15504_320;
  wire  T_15504_321;
  wire  T_15504_322;
  wire  T_15504_323;
  wire  T_15504_324;
  wire  T_15504_325;
  wire  T_15504_326;
  wire  T_15504_327;
  wire  T_15504_328;
  wire  T_15504_329;
  wire  T_15504_330;
  wire  T_15504_331;
  wire  T_15504_332;
  wire  T_15504_333;
  wire  T_15504_334;
  wire  T_15504_335;
  wire  T_15504_336;
  wire  T_15504_337;
  wire  T_15504_338;
  wire  T_15504_339;
  wire  T_15504_340;
  wire  T_15504_341;
  wire  T_15504_342;
  wire  T_15504_343;
  wire  T_15504_344;
  wire  T_15504_345;
  wire  T_15504_346;
  wire  T_15504_347;
  wire  T_15504_348;
  wire  T_15504_349;
  wire  T_15504_350;
  wire  T_15504_351;
  wire  T_15504_352;
  wire  T_15504_353;
  wire  T_15504_354;
  wire  T_15504_355;
  wire  T_15504_356;
  wire  T_15504_357;
  wire  T_15504_358;
  wire  T_15504_359;
  wire  T_15504_360;
  wire  T_15504_361;
  wire  T_15504_362;
  wire  T_15504_363;
  wire  T_15504_364;
  wire  T_15504_365;
  wire  T_15504_366;
  wire  T_15504_367;
  wire  T_15504_368;
  wire  T_15504_369;
  wire  T_15504_370;
  wire  T_15504_371;
  wire  T_15504_372;
  wire  T_15504_373;
  wire  T_15504_374;
  wire  T_15504_375;
  wire  T_15504_376;
  wire  T_15504_377;
  wire  T_15504_378;
  wire  T_15504_379;
  wire  T_15504_380;
  wire  T_15504_381;
  wire  T_15504_382;
  wire  T_15504_383;
  wire  T_15504_384;
  wire  T_15504_385;
  wire  T_15504_386;
  wire  T_15504_387;
  wire  T_15504_388;
  wire  T_15504_389;
  wire  T_15504_390;
  wire  T_15504_391;
  wire  T_15504_392;
  wire  T_15504_393;
  wire  T_15504_394;
  wire  T_15504_395;
  wire  T_15504_396;
  wire  T_15504_397;
  wire  T_15504_398;
  wire  T_15504_399;
  wire  T_15504_400;
  wire  T_15504_401;
  wire  T_15504_402;
  wire  T_15504_403;
  wire  T_15504_404;
  wire  T_15504_405;
  wire  T_15504_406;
  wire  T_15504_407;
  wire  T_15504_408;
  wire  T_15504_409;
  wire  T_15504_410;
  wire  T_15504_411;
  wire  T_15504_412;
  wire  T_15504_413;
  wire  T_15504_414;
  wire  T_15504_415;
  wire  T_15504_416;
  wire  T_15504_417;
  wire  T_15504_418;
  wire  T_15504_419;
  wire  T_15504_420;
  wire  T_15504_421;
  wire  T_15504_422;
  wire  T_15504_423;
  wire  T_15504_424;
  wire  T_15504_425;
  wire  T_15504_426;
  wire  T_15504_427;
  wire  T_15504_428;
  wire  T_15504_429;
  wire  T_15504_430;
  wire  T_15504_431;
  wire  T_15504_432;
  wire  T_15504_433;
  wire  T_15504_434;
  wire  T_15504_435;
  wire  T_15504_436;
  wire  T_15504_437;
  wire  T_15504_438;
  wire  T_15504_439;
  wire  T_15504_440;
  wire  T_15504_441;
  wire  T_15504_442;
  wire  T_15504_443;
  wire  T_15504_444;
  wire  T_15504_445;
  wire  T_15504_446;
  wire  T_15504_447;
  wire  T_15504_448;
  wire  T_15504_449;
  wire  T_15504_450;
  wire  T_15504_451;
  wire  T_15504_452;
  wire  T_15504_453;
  wire  T_15504_454;
  wire  T_15504_455;
  wire  T_15504_456;
  wire  T_15504_457;
  wire  T_15504_458;
  wire  T_15504_459;
  wire  T_15504_460;
  wire  T_15504_461;
  wire  T_15504_462;
  wire  T_15504_463;
  wire  T_15504_464;
  wire  T_15504_465;
  wire  T_15504_466;
  wire  T_15504_467;
  wire  T_15504_468;
  wire  T_15504_469;
  wire  T_15504_470;
  wire  T_15504_471;
  wire  T_15504_472;
  wire  T_15504_473;
  wire  T_15504_474;
  wire  T_15504_475;
  wire  T_15504_476;
  wire  T_15504_477;
  wire  T_15504_478;
  wire  T_15504_479;
  wire  T_15504_480;
  wire  T_15504_481;
  wire  T_15504_482;
  wire  T_15504_483;
  wire  T_15504_484;
  wire  T_15504_485;
  wire  T_15504_486;
  wire  T_15504_487;
  wire  T_15504_488;
  wire  T_15504_489;
  wire  T_15504_490;
  wire  T_15504_491;
  wire  T_15504_492;
  wire  T_15504_493;
  wire  T_15504_494;
  wire  T_15504_495;
  wire  T_15504_496;
  wire  T_15504_497;
  wire  T_15504_498;
  wire  T_15504_499;
  wire  T_15504_500;
  wire  T_15504_501;
  wire  T_15504_502;
  wire  T_15504_503;
  wire  T_15504_504;
  wire  T_15504_505;
  wire  T_15504_506;
  wire  T_15504_507;
  wire  T_15504_508;
  wire  T_15504_509;
  wire  T_15504_510;
  wire  T_15504_511;
  wire  T_16265;
  wire  T_16266;
  wire  T_16267;
  wire  T_16268;
  wire  T_16269;
  wire  T_16270;
  wire  T_16271;
  wire  T_16272;
  wire  T_16273;
  wire  T_16274;
  wire  T_16275;
  wire  T_16276;
  wire  T_16277;
  wire  T_16278;
  wire  T_16279;
  wire  T_16280;
  wire  T_16281;
  wire  T_16282;
  wire  T_16283;
  wire  T_16284;
  wire  T_16285;
  wire  T_16286;
  wire  T_16287;
  wire  T_16288;
  wire  T_16289;
  wire  T_16290;
  wire  T_16291;
  wire  T_16292;
  wire  T_16293;
  wire  T_16294;
  wire  T_16295;
  wire  T_16300;
  wire  T_16301;
  wire  T_16302;
  wire  T_16303;
  wire  T_16304;
  wire  T_16305;
  wire  T_16306;
  wire  T_16307;
  wire  T_16308;
  wire  T_16309;
  wire  T_16310;
  wire  T_16311;
  wire  T_16312;
  wire  T_16313;
  wire  T_16314;
  wire  T_16315;
  wire  T_16316;
  wire  T_16317;
  wire  T_16318;
  wire  T_16509;
  wire  T_16510;
  wire  T_16511;
  wire  T_16512;
  wire  T_16513;
  wire  T_16514;
  wire  T_16515;
  wire  T_16516;
  wire  T_16517;
  wire  T_16518;
  wire  T_16519;
  wire  T_16520;
  wire  T_16521;
  wire  T_16522;
  wire  T_16523;
  wire  T_16524;
  wire  T_16525;
  wire  T_16526;
  wire  T_16527;
  wire  T_16528;
  wire  T_16529;
  wire  T_16530;
  wire  T_16531;
  wire  T_16532;
  wire  T_16533;
  wire  T_16534;
  wire  T_16535;
  wire  T_16536;
  wire  T_16537;
  wire  T_16538;
  wire  T_16539;
  wire  T_16544;
  wire  T_16545;
  wire  T_16546;
  wire  T_16547;
  wire  T_16548;
  wire  T_16549;
  wire  T_16550;
  wire  T_16551;
  wire  T_16552;
  wire  T_16553;
  wire  T_16554;
  wire  T_16555;
  wire  T_16556;
  wire  T_16557;
  wire  T_16558;
  wire  T_16559;
  wire  T_16560;
  wire  T_16561;
  wire  T_16562;
  wire  T_18228_0;
  wire  T_18228_1;
  wire  T_18228_2;
  wire  T_18228_3;
  wire  T_18228_4;
  wire  T_18228_5;
  wire  T_18228_6;
  wire  T_18228_7;
  wire  T_18228_8;
  wire  T_18228_9;
  wire  T_18228_10;
  wire  T_18228_11;
  wire  T_18228_12;
  wire  T_18228_13;
  wire  T_18228_14;
  wire  T_18228_15;
  wire  T_18228_16;
  wire  T_18228_17;
  wire  T_18228_18;
  wire  T_18228_19;
  wire  T_18228_20;
  wire  T_18228_21;
  wire  T_18228_22;
  wire  T_18228_23;
  wire  T_18228_24;
  wire  T_18228_25;
  wire  T_18228_26;
  wire  T_18228_27;
  wire  T_18228_28;
  wire  T_18228_29;
  wire  T_18228_30;
  wire  T_18228_31;
  wire  T_18228_32;
  wire  T_18228_33;
  wire  T_18228_34;
  wire  T_18228_35;
  wire  T_18228_36;
  wire  T_18228_37;
  wire  T_18228_38;
  wire  T_18228_39;
  wire  T_18228_40;
  wire  T_18228_41;
  wire  T_18228_42;
  wire  T_18228_43;
  wire  T_18228_44;
  wire  T_18228_45;
  wire  T_18228_46;
  wire  T_18228_47;
  wire  T_18228_48;
  wire  T_18228_49;
  wire  T_18228_50;
  wire  T_18228_51;
  wire  T_18228_52;
  wire  T_18228_53;
  wire  T_18228_54;
  wire  T_18228_55;
  wire  T_18228_56;
  wire  T_18228_57;
  wire  T_18228_58;
  wire  T_18228_59;
  wire  T_18228_60;
  wire  T_18228_61;
  wire  T_18228_62;
  wire  T_18228_63;
  wire  T_18228_64;
  wire  T_18228_65;
  wire  T_18228_66;
  wire  T_18228_67;
  wire  T_18228_68;
  wire  T_18228_69;
  wire  T_18228_70;
  wire  T_18228_71;
  wire  T_18228_72;
  wire  T_18228_73;
  wire  T_18228_74;
  wire  T_18228_75;
  wire  T_18228_76;
  wire  T_18228_77;
  wire  T_18228_78;
  wire  T_18228_79;
  wire  T_18228_80;
  wire  T_18228_81;
  wire  T_18228_82;
  wire  T_18228_83;
  wire  T_18228_84;
  wire  T_18228_85;
  wire  T_18228_86;
  wire  T_18228_87;
  wire  T_18228_88;
  wire  T_18228_89;
  wire  T_18228_90;
  wire  T_18228_91;
  wire  T_18228_92;
  wire  T_18228_93;
  wire  T_18228_94;
  wire  T_18228_95;
  wire  T_18228_96;
  wire  T_18228_97;
  wire  T_18228_98;
  wire  T_18228_99;
  wire  T_18228_100;
  wire  T_18228_101;
  wire  T_18228_102;
  wire  T_18228_103;
  wire  T_18228_104;
  wire  T_18228_105;
  wire  T_18228_106;
  wire  T_18228_107;
  wire  T_18228_108;
  wire  T_18228_109;
  wire  T_18228_110;
  wire  T_18228_111;
  wire  T_18228_112;
  wire  T_18228_113;
  wire  T_18228_114;
  wire  T_18228_115;
  wire  T_18228_116;
  wire  T_18228_117;
  wire  T_18228_118;
  wire  T_18228_119;
  wire  T_18228_120;
  wire  T_18228_121;
  wire  T_18228_122;
  wire  T_18228_123;
  wire  T_18228_124;
  wire  T_18228_125;
  wire  T_18228_126;
  wire  T_18228_127;
  wire  T_18228_128;
  wire  T_18228_129;
  wire  T_18228_130;
  wire  T_18228_131;
  wire  T_18228_132;
  wire  T_18228_133;
  wire  T_18228_134;
  wire  T_18228_135;
  wire  T_18228_136;
  wire  T_18228_137;
  wire  T_18228_138;
  wire  T_18228_139;
  wire  T_18228_140;
  wire  T_18228_141;
  wire  T_18228_142;
  wire  T_18228_143;
  wire  T_18228_144;
  wire  T_18228_145;
  wire  T_18228_146;
  wire  T_18228_147;
  wire  T_18228_148;
  wire  T_18228_149;
  wire  T_18228_150;
  wire  T_18228_151;
  wire  T_18228_152;
  wire  T_18228_153;
  wire  T_18228_154;
  wire  T_18228_155;
  wire  T_18228_156;
  wire  T_18228_157;
  wire  T_18228_158;
  wire  T_18228_159;
  wire  T_18228_160;
  wire  T_18228_161;
  wire  T_18228_162;
  wire  T_18228_163;
  wire  T_18228_164;
  wire  T_18228_165;
  wire  T_18228_166;
  wire  T_18228_167;
  wire  T_18228_168;
  wire  T_18228_169;
  wire  T_18228_170;
  wire  T_18228_171;
  wire  T_18228_172;
  wire  T_18228_173;
  wire  T_18228_174;
  wire  T_18228_175;
  wire  T_18228_176;
  wire  T_18228_177;
  wire  T_18228_178;
  wire  T_18228_179;
  wire  T_18228_180;
  wire  T_18228_181;
  wire  T_18228_182;
  wire  T_18228_183;
  wire  T_18228_184;
  wire  T_18228_185;
  wire  T_18228_186;
  wire  T_18228_187;
  wire  T_18228_188;
  wire  T_18228_189;
  wire  T_18228_190;
  wire  T_18228_191;
  wire  T_18228_192;
  wire  T_18228_193;
  wire  T_18228_194;
  wire  T_18228_195;
  wire  T_18228_196;
  wire  T_18228_197;
  wire  T_18228_198;
  wire  T_18228_199;
  wire  T_18228_200;
  wire  T_18228_201;
  wire  T_18228_202;
  wire  T_18228_203;
  wire  T_18228_204;
  wire  T_18228_205;
  wire  T_18228_206;
  wire  T_18228_207;
  wire  T_18228_208;
  wire  T_18228_209;
  wire  T_18228_210;
  wire  T_18228_211;
  wire  T_18228_212;
  wire  T_18228_213;
  wire  T_18228_214;
  wire  T_18228_215;
  wire  T_18228_216;
  wire  T_18228_217;
  wire  T_18228_218;
  wire  T_18228_219;
  wire  T_18228_220;
  wire  T_18228_221;
  wire  T_18228_222;
  wire  T_18228_223;
  wire  T_18228_224;
  wire  T_18228_225;
  wire  T_18228_226;
  wire  T_18228_227;
  wire  T_18228_228;
  wire  T_18228_229;
  wire  T_18228_230;
  wire  T_18228_231;
  wire  T_18228_232;
  wire  T_18228_233;
  wire  T_18228_234;
  wire  T_18228_235;
  wire  T_18228_236;
  wire  T_18228_237;
  wire  T_18228_238;
  wire  T_18228_239;
  wire  T_18228_240;
  wire  T_18228_241;
  wire  T_18228_242;
  wire  T_18228_243;
  wire  T_18228_244;
  wire  T_18228_245;
  wire  T_18228_246;
  wire  T_18228_247;
  wire  T_18228_248;
  wire  T_18228_249;
  wire  T_18228_250;
  wire  T_18228_251;
  wire  T_18228_252;
  wire  T_18228_253;
  wire  T_18228_254;
  wire  T_18228_255;
  wire  T_18228_256;
  wire  T_18228_257;
  wire  T_18228_258;
  wire  T_18228_259;
  wire  T_18228_260;
  wire  T_18228_261;
  wire  T_18228_262;
  wire  T_18228_263;
  wire  T_18228_264;
  wire  T_18228_265;
  wire  T_18228_266;
  wire  T_18228_267;
  wire  T_18228_268;
  wire  T_18228_269;
  wire  T_18228_270;
  wire  T_18228_271;
  wire  T_18228_272;
  wire  T_18228_273;
  wire  T_18228_274;
  wire  T_18228_275;
  wire  T_18228_276;
  wire  T_18228_277;
  wire  T_18228_278;
  wire  T_18228_279;
  wire  T_18228_280;
  wire  T_18228_281;
  wire  T_18228_282;
  wire  T_18228_283;
  wire  T_18228_284;
  wire  T_18228_285;
  wire  T_18228_286;
  wire  T_18228_287;
  wire  T_18228_288;
  wire  T_18228_289;
  wire  T_18228_290;
  wire  T_18228_291;
  wire  T_18228_292;
  wire  T_18228_293;
  wire  T_18228_294;
  wire  T_18228_295;
  wire  T_18228_296;
  wire  T_18228_297;
  wire  T_18228_298;
  wire  T_18228_299;
  wire  T_18228_300;
  wire  T_18228_301;
  wire  T_18228_302;
  wire  T_18228_303;
  wire  T_18228_304;
  wire  T_18228_305;
  wire  T_18228_306;
  wire  T_18228_307;
  wire  T_18228_308;
  wire  T_18228_309;
  wire  T_18228_310;
  wire  T_18228_311;
  wire  T_18228_312;
  wire  T_18228_313;
  wire  T_18228_314;
  wire  T_18228_315;
  wire  T_18228_316;
  wire  T_18228_317;
  wire  T_18228_318;
  wire  T_18228_319;
  wire  T_18228_320;
  wire  T_18228_321;
  wire  T_18228_322;
  wire  T_18228_323;
  wire  T_18228_324;
  wire  T_18228_325;
  wire  T_18228_326;
  wire  T_18228_327;
  wire  T_18228_328;
  wire  T_18228_329;
  wire  T_18228_330;
  wire  T_18228_331;
  wire  T_18228_332;
  wire  T_18228_333;
  wire  T_18228_334;
  wire  T_18228_335;
  wire  T_18228_336;
  wire  T_18228_337;
  wire  T_18228_338;
  wire  T_18228_339;
  wire  T_18228_340;
  wire  T_18228_341;
  wire  T_18228_342;
  wire  T_18228_343;
  wire  T_18228_344;
  wire  T_18228_345;
  wire  T_18228_346;
  wire  T_18228_347;
  wire  T_18228_348;
  wire  T_18228_349;
  wire  T_18228_350;
  wire  T_18228_351;
  wire  T_18228_352;
  wire  T_18228_353;
  wire  T_18228_354;
  wire  T_18228_355;
  wire  T_18228_356;
  wire  T_18228_357;
  wire  T_18228_358;
  wire  T_18228_359;
  wire  T_18228_360;
  wire  T_18228_361;
  wire  T_18228_362;
  wire  T_18228_363;
  wire  T_18228_364;
  wire  T_18228_365;
  wire  T_18228_366;
  wire  T_18228_367;
  wire  T_18228_368;
  wire  T_18228_369;
  wire  T_18228_370;
  wire  T_18228_371;
  wire  T_18228_372;
  wire  T_18228_373;
  wire  T_18228_374;
  wire  T_18228_375;
  wire  T_18228_376;
  wire  T_18228_377;
  wire  T_18228_378;
  wire  T_18228_379;
  wire  T_18228_380;
  wire  T_18228_381;
  wire  T_18228_382;
  wire  T_18228_383;
  wire  T_18228_384;
  wire  T_18228_385;
  wire  T_18228_386;
  wire  T_18228_387;
  wire  T_18228_388;
  wire  T_18228_389;
  wire  T_18228_390;
  wire  T_18228_391;
  wire  T_18228_392;
  wire  T_18228_393;
  wire  T_18228_394;
  wire  T_18228_395;
  wire  T_18228_396;
  wire  T_18228_397;
  wire  T_18228_398;
  wire  T_18228_399;
  wire  T_18228_400;
  wire  T_18228_401;
  wire  T_18228_402;
  wire  T_18228_403;
  wire  T_18228_404;
  wire  T_18228_405;
  wire  T_18228_406;
  wire  T_18228_407;
  wire  T_18228_408;
  wire  T_18228_409;
  wire  T_18228_410;
  wire  T_18228_411;
  wire  T_18228_412;
  wire  T_18228_413;
  wire  T_18228_414;
  wire  T_18228_415;
  wire  T_18228_416;
  wire  T_18228_417;
  wire  T_18228_418;
  wire  T_18228_419;
  wire  T_18228_420;
  wire  T_18228_421;
  wire  T_18228_422;
  wire  T_18228_423;
  wire  T_18228_424;
  wire  T_18228_425;
  wire  T_18228_426;
  wire  T_18228_427;
  wire  T_18228_428;
  wire  T_18228_429;
  wire  T_18228_430;
  wire  T_18228_431;
  wire  T_18228_432;
  wire  T_18228_433;
  wire  T_18228_434;
  wire  T_18228_435;
  wire  T_18228_436;
  wire  T_18228_437;
  wire  T_18228_438;
  wire  T_18228_439;
  wire  T_18228_440;
  wire  T_18228_441;
  wire  T_18228_442;
  wire  T_18228_443;
  wire  T_18228_444;
  wire  T_18228_445;
  wire  T_18228_446;
  wire  T_18228_447;
  wire  T_18228_448;
  wire  T_18228_449;
  wire  T_18228_450;
  wire  T_18228_451;
  wire  T_18228_452;
  wire  T_18228_453;
  wire  T_18228_454;
  wire  T_18228_455;
  wire  T_18228_456;
  wire  T_18228_457;
  wire  T_18228_458;
  wire  T_18228_459;
  wire  T_18228_460;
  wire  T_18228_461;
  wire  T_18228_462;
  wire  T_18228_463;
  wire  T_18228_464;
  wire  T_18228_465;
  wire  T_18228_466;
  wire  T_18228_467;
  wire  T_18228_468;
  wire  T_18228_469;
  wire  T_18228_470;
  wire  T_18228_471;
  wire  T_18228_472;
  wire  T_18228_473;
  wire  T_18228_474;
  wire  T_18228_475;
  wire  T_18228_476;
  wire  T_18228_477;
  wire  T_18228_478;
  wire  T_18228_479;
  wire  T_18228_480;
  wire  T_18228_481;
  wire  T_18228_482;
  wire  T_18228_483;
  wire  T_18228_484;
  wire  T_18228_485;
  wire  T_18228_486;
  wire  T_18228_487;
  wire  T_18228_488;
  wire  T_18228_489;
  wire  T_18228_490;
  wire  T_18228_491;
  wire  T_18228_492;
  wire  T_18228_493;
  wire  T_18228_494;
  wire  T_18228_495;
  wire  T_18228_496;
  wire  T_18228_497;
  wire  T_18228_498;
  wire  T_18228_499;
  wire  T_18228_500;
  wire  T_18228_501;
  wire  T_18228_502;
  wire  T_18228_503;
  wire  T_18228_504;
  wire  T_18228_505;
  wire  T_18228_506;
  wire  T_18228_507;
  wire  T_18228_508;
  wire  T_18228_509;
  wire  T_18228_510;
  wire  T_18228_511;
  wire  T_18989;
  wire  T_18990;
  wire  T_18991;
  wire  T_18992;
  wire  T_18993;
  wire  T_18994;
  wire  T_18995;
  wire  T_18996;
  wire  T_18997;
  wire  T_18998;
  wire  T_18999;
  wire  T_19000;
  wire  T_19001;
  wire  T_19002;
  wire  T_19003;
  wire  T_19004;
  wire  T_19005;
  wire  T_19006;
  wire  T_19007;
  wire  T_19008;
  wire  T_19009;
  wire  T_19010;
  wire  T_19011;
  wire  T_19012;
  wire  T_19013;
  wire  T_19014;
  wire  T_19015;
  wire  T_19016;
  wire  T_19017;
  wire  T_19018;
  wire  T_19019;
  wire  T_19024;
  wire  T_19025;
  wire  T_19026;
  wire  T_19027;
  wire  T_19028;
  wire  T_19029;
  wire  T_19030;
  wire  T_19031;
  wire  T_19032;
  wire  T_19033;
  wire  T_19034;
  wire  T_19035;
  wire  T_19036;
  wire  T_19037;
  wire  T_19038;
  wire  T_19039;
  wire  T_19040;
  wire  T_19041;
  wire  T_19042;
  wire  T_19233;
  wire  T_19234;
  wire  T_19235;
  wire  T_19236;
  wire  T_19237;
  wire  T_19238;
  wire  T_19239;
  wire  T_19240;
  wire  T_19241;
  wire  T_19242;
  wire  T_19243;
  wire  T_19244;
  wire  T_19245;
  wire  T_19246;
  wire  T_19247;
  wire  T_19248;
  wire  T_19249;
  wire  T_19250;
  wire  T_19251;
  wire  T_19252;
  wire  T_19253;
  wire  T_19254;
  wire  T_19255;
  wire  T_19256;
  wire  T_19257;
  wire  T_19258;
  wire  T_19259;
  wire  T_19260;
  wire  T_19261;
  wire  T_19262;
  wire  T_19263;
  wire  T_19268;
  wire  T_19269;
  wire  T_19270;
  wire  T_19271;
  wire  T_19272;
  wire  T_19273;
  wire  T_19274;
  wire  T_19275;
  wire  T_19276;
  wire  T_19277;
  wire  T_19278;
  wire  T_19279;
  wire  T_19280;
  wire  T_19281;
  wire  T_19282;
  wire  T_19283;
  wire  T_19284;
  wire  T_19285;
  wire  T_19286;
  wire  T_20952_0;
  wire  T_20952_1;
  wire  T_20952_2;
  wire  T_20952_3;
  wire  T_20952_4;
  wire  T_20952_5;
  wire  T_20952_6;
  wire  T_20952_7;
  wire  T_20952_8;
  wire  T_20952_9;
  wire  T_20952_10;
  wire  T_20952_11;
  wire  T_20952_12;
  wire  T_20952_13;
  wire  T_20952_14;
  wire  T_20952_15;
  wire  T_20952_16;
  wire  T_20952_17;
  wire  T_20952_18;
  wire  T_20952_19;
  wire  T_20952_20;
  wire  T_20952_21;
  wire  T_20952_22;
  wire  T_20952_23;
  wire  T_20952_24;
  wire  T_20952_25;
  wire  T_20952_26;
  wire  T_20952_27;
  wire  T_20952_28;
  wire  T_20952_29;
  wire  T_20952_30;
  wire  T_20952_31;
  wire  T_20952_32;
  wire  T_20952_33;
  wire  T_20952_34;
  wire  T_20952_35;
  wire  T_20952_36;
  wire  T_20952_37;
  wire  T_20952_38;
  wire  T_20952_39;
  wire  T_20952_40;
  wire  T_20952_41;
  wire  T_20952_42;
  wire  T_20952_43;
  wire  T_20952_44;
  wire  T_20952_45;
  wire  T_20952_46;
  wire  T_20952_47;
  wire  T_20952_48;
  wire  T_20952_49;
  wire  T_20952_50;
  wire  T_20952_51;
  wire  T_20952_52;
  wire  T_20952_53;
  wire  T_20952_54;
  wire  T_20952_55;
  wire  T_20952_56;
  wire  T_20952_57;
  wire  T_20952_58;
  wire  T_20952_59;
  wire  T_20952_60;
  wire  T_20952_61;
  wire  T_20952_62;
  wire  T_20952_63;
  wire  T_20952_64;
  wire  T_20952_65;
  wire  T_20952_66;
  wire  T_20952_67;
  wire  T_20952_68;
  wire  T_20952_69;
  wire  T_20952_70;
  wire  T_20952_71;
  wire  T_20952_72;
  wire  T_20952_73;
  wire  T_20952_74;
  wire  T_20952_75;
  wire  T_20952_76;
  wire  T_20952_77;
  wire  T_20952_78;
  wire  T_20952_79;
  wire  T_20952_80;
  wire  T_20952_81;
  wire  T_20952_82;
  wire  T_20952_83;
  wire  T_20952_84;
  wire  T_20952_85;
  wire  T_20952_86;
  wire  T_20952_87;
  wire  T_20952_88;
  wire  T_20952_89;
  wire  T_20952_90;
  wire  T_20952_91;
  wire  T_20952_92;
  wire  T_20952_93;
  wire  T_20952_94;
  wire  T_20952_95;
  wire  T_20952_96;
  wire  T_20952_97;
  wire  T_20952_98;
  wire  T_20952_99;
  wire  T_20952_100;
  wire  T_20952_101;
  wire  T_20952_102;
  wire  T_20952_103;
  wire  T_20952_104;
  wire  T_20952_105;
  wire  T_20952_106;
  wire  T_20952_107;
  wire  T_20952_108;
  wire  T_20952_109;
  wire  T_20952_110;
  wire  T_20952_111;
  wire  T_20952_112;
  wire  T_20952_113;
  wire  T_20952_114;
  wire  T_20952_115;
  wire  T_20952_116;
  wire  T_20952_117;
  wire  T_20952_118;
  wire  T_20952_119;
  wire  T_20952_120;
  wire  T_20952_121;
  wire  T_20952_122;
  wire  T_20952_123;
  wire  T_20952_124;
  wire  T_20952_125;
  wire  T_20952_126;
  wire  T_20952_127;
  wire  T_20952_128;
  wire  T_20952_129;
  wire  T_20952_130;
  wire  T_20952_131;
  wire  T_20952_132;
  wire  T_20952_133;
  wire  T_20952_134;
  wire  T_20952_135;
  wire  T_20952_136;
  wire  T_20952_137;
  wire  T_20952_138;
  wire  T_20952_139;
  wire  T_20952_140;
  wire  T_20952_141;
  wire  T_20952_142;
  wire  T_20952_143;
  wire  T_20952_144;
  wire  T_20952_145;
  wire  T_20952_146;
  wire  T_20952_147;
  wire  T_20952_148;
  wire  T_20952_149;
  wire  T_20952_150;
  wire  T_20952_151;
  wire  T_20952_152;
  wire  T_20952_153;
  wire  T_20952_154;
  wire  T_20952_155;
  wire  T_20952_156;
  wire  T_20952_157;
  wire  T_20952_158;
  wire  T_20952_159;
  wire  T_20952_160;
  wire  T_20952_161;
  wire  T_20952_162;
  wire  T_20952_163;
  wire  T_20952_164;
  wire  T_20952_165;
  wire  T_20952_166;
  wire  T_20952_167;
  wire  T_20952_168;
  wire  T_20952_169;
  wire  T_20952_170;
  wire  T_20952_171;
  wire  T_20952_172;
  wire  T_20952_173;
  wire  T_20952_174;
  wire  T_20952_175;
  wire  T_20952_176;
  wire  T_20952_177;
  wire  T_20952_178;
  wire  T_20952_179;
  wire  T_20952_180;
  wire  T_20952_181;
  wire  T_20952_182;
  wire  T_20952_183;
  wire  T_20952_184;
  wire  T_20952_185;
  wire  T_20952_186;
  wire  T_20952_187;
  wire  T_20952_188;
  wire  T_20952_189;
  wire  T_20952_190;
  wire  T_20952_191;
  wire  T_20952_192;
  wire  T_20952_193;
  wire  T_20952_194;
  wire  T_20952_195;
  wire  T_20952_196;
  wire  T_20952_197;
  wire  T_20952_198;
  wire  T_20952_199;
  wire  T_20952_200;
  wire  T_20952_201;
  wire  T_20952_202;
  wire  T_20952_203;
  wire  T_20952_204;
  wire  T_20952_205;
  wire  T_20952_206;
  wire  T_20952_207;
  wire  T_20952_208;
  wire  T_20952_209;
  wire  T_20952_210;
  wire  T_20952_211;
  wire  T_20952_212;
  wire  T_20952_213;
  wire  T_20952_214;
  wire  T_20952_215;
  wire  T_20952_216;
  wire  T_20952_217;
  wire  T_20952_218;
  wire  T_20952_219;
  wire  T_20952_220;
  wire  T_20952_221;
  wire  T_20952_222;
  wire  T_20952_223;
  wire  T_20952_224;
  wire  T_20952_225;
  wire  T_20952_226;
  wire  T_20952_227;
  wire  T_20952_228;
  wire  T_20952_229;
  wire  T_20952_230;
  wire  T_20952_231;
  wire  T_20952_232;
  wire  T_20952_233;
  wire  T_20952_234;
  wire  T_20952_235;
  wire  T_20952_236;
  wire  T_20952_237;
  wire  T_20952_238;
  wire  T_20952_239;
  wire  T_20952_240;
  wire  T_20952_241;
  wire  T_20952_242;
  wire  T_20952_243;
  wire  T_20952_244;
  wire  T_20952_245;
  wire  T_20952_246;
  wire  T_20952_247;
  wire  T_20952_248;
  wire  T_20952_249;
  wire  T_20952_250;
  wire  T_20952_251;
  wire  T_20952_252;
  wire  T_20952_253;
  wire  T_20952_254;
  wire  T_20952_255;
  wire  T_20952_256;
  wire  T_20952_257;
  wire  T_20952_258;
  wire  T_20952_259;
  wire  T_20952_260;
  wire  T_20952_261;
  wire  T_20952_262;
  wire  T_20952_263;
  wire  T_20952_264;
  wire  T_20952_265;
  wire  T_20952_266;
  wire  T_20952_267;
  wire  T_20952_268;
  wire  T_20952_269;
  wire  T_20952_270;
  wire  T_20952_271;
  wire  T_20952_272;
  wire  T_20952_273;
  wire  T_20952_274;
  wire  T_20952_275;
  wire  T_20952_276;
  wire  T_20952_277;
  wire  T_20952_278;
  wire  T_20952_279;
  wire  T_20952_280;
  wire  T_20952_281;
  wire  T_20952_282;
  wire  T_20952_283;
  wire  T_20952_284;
  wire  T_20952_285;
  wire  T_20952_286;
  wire  T_20952_287;
  wire  T_20952_288;
  wire  T_20952_289;
  wire  T_20952_290;
  wire  T_20952_291;
  wire  T_20952_292;
  wire  T_20952_293;
  wire  T_20952_294;
  wire  T_20952_295;
  wire  T_20952_296;
  wire  T_20952_297;
  wire  T_20952_298;
  wire  T_20952_299;
  wire  T_20952_300;
  wire  T_20952_301;
  wire  T_20952_302;
  wire  T_20952_303;
  wire  T_20952_304;
  wire  T_20952_305;
  wire  T_20952_306;
  wire  T_20952_307;
  wire  T_20952_308;
  wire  T_20952_309;
  wire  T_20952_310;
  wire  T_20952_311;
  wire  T_20952_312;
  wire  T_20952_313;
  wire  T_20952_314;
  wire  T_20952_315;
  wire  T_20952_316;
  wire  T_20952_317;
  wire  T_20952_318;
  wire  T_20952_319;
  wire  T_20952_320;
  wire  T_20952_321;
  wire  T_20952_322;
  wire  T_20952_323;
  wire  T_20952_324;
  wire  T_20952_325;
  wire  T_20952_326;
  wire  T_20952_327;
  wire  T_20952_328;
  wire  T_20952_329;
  wire  T_20952_330;
  wire  T_20952_331;
  wire  T_20952_332;
  wire  T_20952_333;
  wire  T_20952_334;
  wire  T_20952_335;
  wire  T_20952_336;
  wire  T_20952_337;
  wire  T_20952_338;
  wire  T_20952_339;
  wire  T_20952_340;
  wire  T_20952_341;
  wire  T_20952_342;
  wire  T_20952_343;
  wire  T_20952_344;
  wire  T_20952_345;
  wire  T_20952_346;
  wire  T_20952_347;
  wire  T_20952_348;
  wire  T_20952_349;
  wire  T_20952_350;
  wire  T_20952_351;
  wire  T_20952_352;
  wire  T_20952_353;
  wire  T_20952_354;
  wire  T_20952_355;
  wire  T_20952_356;
  wire  T_20952_357;
  wire  T_20952_358;
  wire  T_20952_359;
  wire  T_20952_360;
  wire  T_20952_361;
  wire  T_20952_362;
  wire  T_20952_363;
  wire  T_20952_364;
  wire  T_20952_365;
  wire  T_20952_366;
  wire  T_20952_367;
  wire  T_20952_368;
  wire  T_20952_369;
  wire  T_20952_370;
  wire  T_20952_371;
  wire  T_20952_372;
  wire  T_20952_373;
  wire  T_20952_374;
  wire  T_20952_375;
  wire  T_20952_376;
  wire  T_20952_377;
  wire  T_20952_378;
  wire  T_20952_379;
  wire  T_20952_380;
  wire  T_20952_381;
  wire  T_20952_382;
  wire  T_20952_383;
  wire  T_20952_384;
  wire  T_20952_385;
  wire  T_20952_386;
  wire  T_20952_387;
  wire  T_20952_388;
  wire  T_20952_389;
  wire  T_20952_390;
  wire  T_20952_391;
  wire  T_20952_392;
  wire  T_20952_393;
  wire  T_20952_394;
  wire  T_20952_395;
  wire  T_20952_396;
  wire  T_20952_397;
  wire  T_20952_398;
  wire  T_20952_399;
  wire  T_20952_400;
  wire  T_20952_401;
  wire  T_20952_402;
  wire  T_20952_403;
  wire  T_20952_404;
  wire  T_20952_405;
  wire  T_20952_406;
  wire  T_20952_407;
  wire  T_20952_408;
  wire  T_20952_409;
  wire  T_20952_410;
  wire  T_20952_411;
  wire  T_20952_412;
  wire  T_20952_413;
  wire  T_20952_414;
  wire  T_20952_415;
  wire  T_20952_416;
  wire  T_20952_417;
  wire  T_20952_418;
  wire  T_20952_419;
  wire  T_20952_420;
  wire  T_20952_421;
  wire  T_20952_422;
  wire  T_20952_423;
  wire  T_20952_424;
  wire  T_20952_425;
  wire  T_20952_426;
  wire  T_20952_427;
  wire  T_20952_428;
  wire  T_20952_429;
  wire  T_20952_430;
  wire  T_20952_431;
  wire  T_20952_432;
  wire  T_20952_433;
  wire  T_20952_434;
  wire  T_20952_435;
  wire  T_20952_436;
  wire  T_20952_437;
  wire  T_20952_438;
  wire  T_20952_439;
  wire  T_20952_440;
  wire  T_20952_441;
  wire  T_20952_442;
  wire  T_20952_443;
  wire  T_20952_444;
  wire  T_20952_445;
  wire  T_20952_446;
  wire  T_20952_447;
  wire  T_20952_448;
  wire  T_20952_449;
  wire  T_20952_450;
  wire  T_20952_451;
  wire  T_20952_452;
  wire  T_20952_453;
  wire  T_20952_454;
  wire  T_20952_455;
  wire  T_20952_456;
  wire  T_20952_457;
  wire  T_20952_458;
  wire  T_20952_459;
  wire  T_20952_460;
  wire  T_20952_461;
  wire  T_20952_462;
  wire  T_20952_463;
  wire  T_20952_464;
  wire  T_20952_465;
  wire  T_20952_466;
  wire  T_20952_467;
  wire  T_20952_468;
  wire  T_20952_469;
  wire  T_20952_470;
  wire  T_20952_471;
  wire  T_20952_472;
  wire  T_20952_473;
  wire  T_20952_474;
  wire  T_20952_475;
  wire  T_20952_476;
  wire  T_20952_477;
  wire  T_20952_478;
  wire  T_20952_479;
  wire  T_20952_480;
  wire  T_20952_481;
  wire  T_20952_482;
  wire  T_20952_483;
  wire  T_20952_484;
  wire  T_20952_485;
  wire  T_20952_486;
  wire  T_20952_487;
  wire  T_20952_488;
  wire  T_20952_489;
  wire  T_20952_490;
  wire  T_20952_491;
  wire  T_20952_492;
  wire  T_20952_493;
  wire  T_20952_494;
  wire  T_20952_495;
  wire  T_20952_496;
  wire  T_20952_497;
  wire  T_20952_498;
  wire  T_20952_499;
  wire  T_20952_500;
  wire  T_20952_501;
  wire  T_20952_502;
  wire  T_20952_503;
  wire  T_20952_504;
  wire  T_20952_505;
  wire  T_20952_506;
  wire  T_20952_507;
  wire  T_20952_508;
  wire  T_20952_509;
  wire  T_20952_510;
  wire  T_20952_511;
  wire  T_21713;
  wire  T_21714;
  wire  T_21715;
  wire  T_21716;
  wire  T_21717;
  wire  T_21718;
  wire  T_21719;
  wire  T_21720;
  wire  T_21721;
  wire  T_21722;
  wire  T_21723;
  wire  T_21724;
  wire  T_21725;
  wire  T_21726;
  wire  T_21727;
  wire  T_21728;
  wire  T_21729;
  wire  T_21730;
  wire  T_21731;
  wire  T_21732;
  wire  T_21733;
  wire  T_21734;
  wire  T_21735;
  wire  T_21736;
  wire  T_21737;
  wire  T_21738;
  wire  T_21739;
  wire  T_21740;
  wire  T_21741;
  wire  T_21742;
  wire  T_21743;
  wire  T_21748;
  wire  T_21749;
  wire  T_21750;
  wire  T_21751;
  wire  T_21752;
  wire  T_21753;
  wire  T_21754;
  wire  T_21755;
  wire  T_21756;
  wire  T_21757;
  wire  T_21758;
  wire  T_21759;
  wire  T_21760;
  wire  T_21761;
  wire  T_21762;
  wire  T_21763;
  wire  T_21764;
  wire  T_21765;
  wire  T_21766;
  wire  T_21957;
  wire  T_21958;
  wire  T_21959;
  wire  T_21960;
  wire  T_21961;
  wire  T_21962;
  wire  T_21963;
  wire  T_21964;
  wire  T_21965;
  wire  T_21966;
  wire  T_21967;
  wire  T_21968;
  wire  T_21969;
  wire  T_21970;
  wire  T_21971;
  wire  T_21972;
  wire  T_21973;
  wire  T_21974;
  wire  T_21975;
  wire  T_21976;
  wire  T_21977;
  wire  T_21978;
  wire  T_21979;
  wire  T_21980;
  wire  T_21981;
  wire  T_21982;
  wire  T_21983;
  wire  T_21984;
  wire  T_21985;
  wire  T_21986;
  wire  T_21987;
  wire  T_21992;
  wire  T_21993;
  wire  T_21994;
  wire  T_21995;
  wire  T_21996;
  wire  T_21997;
  wire  T_21998;
  wire  T_21999;
  wire  T_22000;
  wire  T_22001;
  wire  T_22002;
  wire  T_22003;
  wire  T_22004;
  wire  T_22005;
  wire  T_22006;
  wire  T_22007;
  wire  T_22008;
  wire  T_22009;
  wire  T_22010;
  wire  T_23676_0;
  wire  T_23676_1;
  wire  T_23676_2;
  wire  T_23676_3;
  wire  T_23676_4;
  wire  T_23676_5;
  wire  T_23676_6;
  wire  T_23676_7;
  wire  T_23676_8;
  wire  T_23676_9;
  wire  T_23676_10;
  wire  T_23676_11;
  wire  T_23676_12;
  wire  T_23676_13;
  wire  T_23676_14;
  wire  T_23676_15;
  wire  T_23676_16;
  wire  T_23676_17;
  wire  T_23676_18;
  wire  T_23676_19;
  wire  T_23676_20;
  wire  T_23676_21;
  wire  T_23676_22;
  wire  T_23676_23;
  wire  T_23676_24;
  wire  T_23676_25;
  wire  T_23676_26;
  wire  T_23676_27;
  wire  T_23676_28;
  wire  T_23676_29;
  wire  T_23676_30;
  wire  T_23676_31;
  wire  T_23676_32;
  wire  T_23676_33;
  wire  T_23676_34;
  wire  T_23676_35;
  wire  T_23676_36;
  wire  T_23676_37;
  wire  T_23676_38;
  wire  T_23676_39;
  wire  T_23676_40;
  wire  T_23676_41;
  wire  T_23676_42;
  wire  T_23676_43;
  wire  T_23676_44;
  wire  T_23676_45;
  wire  T_23676_46;
  wire  T_23676_47;
  wire  T_23676_48;
  wire  T_23676_49;
  wire  T_23676_50;
  wire  T_23676_51;
  wire  T_23676_52;
  wire  T_23676_53;
  wire  T_23676_54;
  wire  T_23676_55;
  wire  T_23676_56;
  wire  T_23676_57;
  wire  T_23676_58;
  wire  T_23676_59;
  wire  T_23676_60;
  wire  T_23676_61;
  wire  T_23676_62;
  wire  T_23676_63;
  wire  T_23676_64;
  wire  T_23676_65;
  wire  T_23676_66;
  wire  T_23676_67;
  wire  T_23676_68;
  wire  T_23676_69;
  wire  T_23676_70;
  wire  T_23676_71;
  wire  T_23676_72;
  wire  T_23676_73;
  wire  T_23676_74;
  wire  T_23676_75;
  wire  T_23676_76;
  wire  T_23676_77;
  wire  T_23676_78;
  wire  T_23676_79;
  wire  T_23676_80;
  wire  T_23676_81;
  wire  T_23676_82;
  wire  T_23676_83;
  wire  T_23676_84;
  wire  T_23676_85;
  wire  T_23676_86;
  wire  T_23676_87;
  wire  T_23676_88;
  wire  T_23676_89;
  wire  T_23676_90;
  wire  T_23676_91;
  wire  T_23676_92;
  wire  T_23676_93;
  wire  T_23676_94;
  wire  T_23676_95;
  wire  T_23676_96;
  wire  T_23676_97;
  wire  T_23676_98;
  wire  T_23676_99;
  wire  T_23676_100;
  wire  T_23676_101;
  wire  T_23676_102;
  wire  T_23676_103;
  wire  T_23676_104;
  wire  T_23676_105;
  wire  T_23676_106;
  wire  T_23676_107;
  wire  T_23676_108;
  wire  T_23676_109;
  wire  T_23676_110;
  wire  T_23676_111;
  wire  T_23676_112;
  wire  T_23676_113;
  wire  T_23676_114;
  wire  T_23676_115;
  wire  T_23676_116;
  wire  T_23676_117;
  wire  T_23676_118;
  wire  T_23676_119;
  wire  T_23676_120;
  wire  T_23676_121;
  wire  T_23676_122;
  wire  T_23676_123;
  wire  T_23676_124;
  wire  T_23676_125;
  wire  T_23676_126;
  wire  T_23676_127;
  wire  T_23676_128;
  wire  T_23676_129;
  wire  T_23676_130;
  wire  T_23676_131;
  wire  T_23676_132;
  wire  T_23676_133;
  wire  T_23676_134;
  wire  T_23676_135;
  wire  T_23676_136;
  wire  T_23676_137;
  wire  T_23676_138;
  wire  T_23676_139;
  wire  T_23676_140;
  wire  T_23676_141;
  wire  T_23676_142;
  wire  T_23676_143;
  wire  T_23676_144;
  wire  T_23676_145;
  wire  T_23676_146;
  wire  T_23676_147;
  wire  T_23676_148;
  wire  T_23676_149;
  wire  T_23676_150;
  wire  T_23676_151;
  wire  T_23676_152;
  wire  T_23676_153;
  wire  T_23676_154;
  wire  T_23676_155;
  wire  T_23676_156;
  wire  T_23676_157;
  wire  T_23676_158;
  wire  T_23676_159;
  wire  T_23676_160;
  wire  T_23676_161;
  wire  T_23676_162;
  wire  T_23676_163;
  wire  T_23676_164;
  wire  T_23676_165;
  wire  T_23676_166;
  wire  T_23676_167;
  wire  T_23676_168;
  wire  T_23676_169;
  wire  T_23676_170;
  wire  T_23676_171;
  wire  T_23676_172;
  wire  T_23676_173;
  wire  T_23676_174;
  wire  T_23676_175;
  wire  T_23676_176;
  wire  T_23676_177;
  wire  T_23676_178;
  wire  T_23676_179;
  wire  T_23676_180;
  wire  T_23676_181;
  wire  T_23676_182;
  wire  T_23676_183;
  wire  T_23676_184;
  wire  T_23676_185;
  wire  T_23676_186;
  wire  T_23676_187;
  wire  T_23676_188;
  wire  T_23676_189;
  wire  T_23676_190;
  wire  T_23676_191;
  wire  T_23676_192;
  wire  T_23676_193;
  wire  T_23676_194;
  wire  T_23676_195;
  wire  T_23676_196;
  wire  T_23676_197;
  wire  T_23676_198;
  wire  T_23676_199;
  wire  T_23676_200;
  wire  T_23676_201;
  wire  T_23676_202;
  wire  T_23676_203;
  wire  T_23676_204;
  wire  T_23676_205;
  wire  T_23676_206;
  wire  T_23676_207;
  wire  T_23676_208;
  wire  T_23676_209;
  wire  T_23676_210;
  wire  T_23676_211;
  wire  T_23676_212;
  wire  T_23676_213;
  wire  T_23676_214;
  wire  T_23676_215;
  wire  T_23676_216;
  wire  T_23676_217;
  wire  T_23676_218;
  wire  T_23676_219;
  wire  T_23676_220;
  wire  T_23676_221;
  wire  T_23676_222;
  wire  T_23676_223;
  wire  T_23676_224;
  wire  T_23676_225;
  wire  T_23676_226;
  wire  T_23676_227;
  wire  T_23676_228;
  wire  T_23676_229;
  wire  T_23676_230;
  wire  T_23676_231;
  wire  T_23676_232;
  wire  T_23676_233;
  wire  T_23676_234;
  wire  T_23676_235;
  wire  T_23676_236;
  wire  T_23676_237;
  wire  T_23676_238;
  wire  T_23676_239;
  wire  T_23676_240;
  wire  T_23676_241;
  wire  T_23676_242;
  wire  T_23676_243;
  wire  T_23676_244;
  wire  T_23676_245;
  wire  T_23676_246;
  wire  T_23676_247;
  wire  T_23676_248;
  wire  T_23676_249;
  wire  T_23676_250;
  wire  T_23676_251;
  wire  T_23676_252;
  wire  T_23676_253;
  wire  T_23676_254;
  wire  T_23676_255;
  wire  T_23676_256;
  wire  T_23676_257;
  wire  T_23676_258;
  wire  T_23676_259;
  wire  T_23676_260;
  wire  T_23676_261;
  wire  T_23676_262;
  wire  T_23676_263;
  wire  T_23676_264;
  wire  T_23676_265;
  wire  T_23676_266;
  wire  T_23676_267;
  wire  T_23676_268;
  wire  T_23676_269;
  wire  T_23676_270;
  wire  T_23676_271;
  wire  T_23676_272;
  wire  T_23676_273;
  wire  T_23676_274;
  wire  T_23676_275;
  wire  T_23676_276;
  wire  T_23676_277;
  wire  T_23676_278;
  wire  T_23676_279;
  wire  T_23676_280;
  wire  T_23676_281;
  wire  T_23676_282;
  wire  T_23676_283;
  wire  T_23676_284;
  wire  T_23676_285;
  wire  T_23676_286;
  wire  T_23676_287;
  wire  T_23676_288;
  wire  T_23676_289;
  wire  T_23676_290;
  wire  T_23676_291;
  wire  T_23676_292;
  wire  T_23676_293;
  wire  T_23676_294;
  wire  T_23676_295;
  wire  T_23676_296;
  wire  T_23676_297;
  wire  T_23676_298;
  wire  T_23676_299;
  wire  T_23676_300;
  wire  T_23676_301;
  wire  T_23676_302;
  wire  T_23676_303;
  wire  T_23676_304;
  wire  T_23676_305;
  wire  T_23676_306;
  wire  T_23676_307;
  wire  T_23676_308;
  wire  T_23676_309;
  wire  T_23676_310;
  wire  T_23676_311;
  wire  T_23676_312;
  wire  T_23676_313;
  wire  T_23676_314;
  wire  T_23676_315;
  wire  T_23676_316;
  wire  T_23676_317;
  wire  T_23676_318;
  wire  T_23676_319;
  wire  T_23676_320;
  wire  T_23676_321;
  wire  T_23676_322;
  wire  T_23676_323;
  wire  T_23676_324;
  wire  T_23676_325;
  wire  T_23676_326;
  wire  T_23676_327;
  wire  T_23676_328;
  wire  T_23676_329;
  wire  T_23676_330;
  wire  T_23676_331;
  wire  T_23676_332;
  wire  T_23676_333;
  wire  T_23676_334;
  wire  T_23676_335;
  wire  T_23676_336;
  wire  T_23676_337;
  wire  T_23676_338;
  wire  T_23676_339;
  wire  T_23676_340;
  wire  T_23676_341;
  wire  T_23676_342;
  wire  T_23676_343;
  wire  T_23676_344;
  wire  T_23676_345;
  wire  T_23676_346;
  wire  T_23676_347;
  wire  T_23676_348;
  wire  T_23676_349;
  wire  T_23676_350;
  wire  T_23676_351;
  wire  T_23676_352;
  wire  T_23676_353;
  wire  T_23676_354;
  wire  T_23676_355;
  wire  T_23676_356;
  wire  T_23676_357;
  wire  T_23676_358;
  wire  T_23676_359;
  wire  T_23676_360;
  wire  T_23676_361;
  wire  T_23676_362;
  wire  T_23676_363;
  wire  T_23676_364;
  wire  T_23676_365;
  wire  T_23676_366;
  wire  T_23676_367;
  wire  T_23676_368;
  wire  T_23676_369;
  wire  T_23676_370;
  wire  T_23676_371;
  wire  T_23676_372;
  wire  T_23676_373;
  wire  T_23676_374;
  wire  T_23676_375;
  wire  T_23676_376;
  wire  T_23676_377;
  wire  T_23676_378;
  wire  T_23676_379;
  wire  T_23676_380;
  wire  T_23676_381;
  wire  T_23676_382;
  wire  T_23676_383;
  wire  T_23676_384;
  wire  T_23676_385;
  wire  T_23676_386;
  wire  T_23676_387;
  wire  T_23676_388;
  wire  T_23676_389;
  wire  T_23676_390;
  wire  T_23676_391;
  wire  T_23676_392;
  wire  T_23676_393;
  wire  T_23676_394;
  wire  T_23676_395;
  wire  T_23676_396;
  wire  T_23676_397;
  wire  T_23676_398;
  wire  T_23676_399;
  wire  T_23676_400;
  wire  T_23676_401;
  wire  T_23676_402;
  wire  T_23676_403;
  wire  T_23676_404;
  wire  T_23676_405;
  wire  T_23676_406;
  wire  T_23676_407;
  wire  T_23676_408;
  wire  T_23676_409;
  wire  T_23676_410;
  wire  T_23676_411;
  wire  T_23676_412;
  wire  T_23676_413;
  wire  T_23676_414;
  wire  T_23676_415;
  wire  T_23676_416;
  wire  T_23676_417;
  wire  T_23676_418;
  wire  T_23676_419;
  wire  T_23676_420;
  wire  T_23676_421;
  wire  T_23676_422;
  wire  T_23676_423;
  wire  T_23676_424;
  wire  T_23676_425;
  wire  T_23676_426;
  wire  T_23676_427;
  wire  T_23676_428;
  wire  T_23676_429;
  wire  T_23676_430;
  wire  T_23676_431;
  wire  T_23676_432;
  wire  T_23676_433;
  wire  T_23676_434;
  wire  T_23676_435;
  wire  T_23676_436;
  wire  T_23676_437;
  wire  T_23676_438;
  wire  T_23676_439;
  wire  T_23676_440;
  wire  T_23676_441;
  wire  T_23676_442;
  wire  T_23676_443;
  wire  T_23676_444;
  wire  T_23676_445;
  wire  T_23676_446;
  wire  T_23676_447;
  wire  T_23676_448;
  wire  T_23676_449;
  wire  T_23676_450;
  wire  T_23676_451;
  wire  T_23676_452;
  wire  T_23676_453;
  wire  T_23676_454;
  wire  T_23676_455;
  wire  T_23676_456;
  wire  T_23676_457;
  wire  T_23676_458;
  wire  T_23676_459;
  wire  T_23676_460;
  wire  T_23676_461;
  wire  T_23676_462;
  wire  T_23676_463;
  wire  T_23676_464;
  wire  T_23676_465;
  wire  T_23676_466;
  wire  T_23676_467;
  wire  T_23676_468;
  wire  T_23676_469;
  wire  T_23676_470;
  wire  T_23676_471;
  wire  T_23676_472;
  wire  T_23676_473;
  wire  T_23676_474;
  wire  T_23676_475;
  wire  T_23676_476;
  wire  T_23676_477;
  wire  T_23676_478;
  wire  T_23676_479;
  wire  T_23676_480;
  wire  T_23676_481;
  wire  T_23676_482;
  wire  T_23676_483;
  wire  T_23676_484;
  wire  T_23676_485;
  wire  T_23676_486;
  wire  T_23676_487;
  wire  T_23676_488;
  wire  T_23676_489;
  wire  T_23676_490;
  wire  T_23676_491;
  wire  T_23676_492;
  wire  T_23676_493;
  wire  T_23676_494;
  wire  T_23676_495;
  wire  T_23676_496;
  wire  T_23676_497;
  wire  T_23676_498;
  wire  T_23676_499;
  wire  T_23676_500;
  wire  T_23676_501;
  wire  T_23676_502;
  wire  T_23676_503;
  wire  T_23676_504;
  wire  T_23676_505;
  wire  T_23676_506;
  wire  T_23676_507;
  wire  T_23676_508;
  wire  T_23676_509;
  wire  T_23676_510;
  wire  T_23676_511;
  wire  T_24191;
  wire  T_24192;
  wire  T_24193;
  wire  T_24194;
  wire  T_24195;
  wire  T_24196;
  wire  T_24201;
  wire  T_24202;
  wire  T_24210;
  wire [1:0] T_24215;
  wire [1:0] T_24216;
  wire [3:0] T_24217;
  wire [1:0] T_24218;
  wire [1:0] T_24219;
  wire [2:0] T_24220;
  wire [4:0] T_24221;
  wire [8:0] T_24222;
  wire  GEN_3;
  wire  GEN_423;
  wire  GEN_424;
  wire  GEN_425;
  wire  GEN_426;
  wire  GEN_427;
  wire  GEN_428;
  wire  GEN_429;
  wire  GEN_430;
  wire  GEN_431;
  wire  GEN_432;
  wire  GEN_433;
  wire  GEN_434;
  wire  GEN_435;
  wire  GEN_436;
  wire  GEN_437;
  wire  GEN_438;
  wire  GEN_439;
  wire  GEN_440;
  wire  GEN_441;
  wire  GEN_442;
  wire  GEN_443;
  wire  GEN_444;
  wire  GEN_445;
  wire  GEN_446;
  wire  GEN_447;
  wire  GEN_448;
  wire  GEN_449;
  wire  GEN_450;
  wire  GEN_451;
  wire  GEN_452;
  wire  GEN_453;
  wire  GEN_454;
  wire  GEN_455;
  wire  GEN_456;
  wire  GEN_457;
  wire  GEN_458;
  wire  GEN_459;
  wire  GEN_460;
  wire  GEN_461;
  wire  GEN_462;
  wire  GEN_463;
  wire  GEN_464;
  wire  GEN_465;
  wire  GEN_466;
  wire  GEN_467;
  wire  GEN_468;
  wire  GEN_469;
  wire  GEN_470;
  wire  GEN_471;
  wire  GEN_472;
  wire  GEN_473;
  wire  GEN_474;
  wire  GEN_475;
  wire  GEN_476;
  wire  GEN_477;
  wire  GEN_478;
  wire  GEN_479;
  wire  GEN_480;
  wire  GEN_481;
  wire  GEN_482;
  wire  GEN_483;
  wire  GEN_484;
  wire  GEN_485;
  wire  GEN_486;
  wire  GEN_487;
  wire  GEN_488;
  wire  GEN_489;
  wire  GEN_490;
  wire  GEN_491;
  wire  GEN_492;
  wire  GEN_493;
  wire  GEN_494;
  wire  GEN_495;
  wire  GEN_496;
  wire  GEN_497;
  wire  GEN_498;
  wire  GEN_499;
  wire  GEN_500;
  wire  GEN_501;
  wire  GEN_502;
  wire  GEN_503;
  wire  GEN_504;
  wire  GEN_505;
  wire  GEN_506;
  wire  GEN_507;
  wire  GEN_508;
  wire  GEN_509;
  wire  GEN_510;
  wire  GEN_511;
  wire  GEN_512;
  wire  GEN_513;
  wire  GEN_514;
  wire  GEN_515;
  wire  GEN_516;
  wire  GEN_517;
  wire  GEN_518;
  wire  GEN_519;
  wire  GEN_520;
  wire  GEN_521;
  wire  GEN_522;
  wire  GEN_523;
  wire  GEN_524;
  wire  GEN_525;
  wire  GEN_526;
  wire  GEN_527;
  wire  GEN_528;
  wire  GEN_529;
  wire  GEN_530;
  wire  GEN_531;
  wire  GEN_532;
  wire  GEN_533;
  wire  GEN_534;
  wire  GEN_535;
  wire  GEN_536;
  wire  GEN_537;
  wire  GEN_538;
  wire  GEN_539;
  wire  GEN_540;
  wire  GEN_541;
  wire  GEN_542;
  wire  GEN_543;
  wire  GEN_544;
  wire  GEN_545;
  wire  GEN_546;
  wire  GEN_547;
  wire  GEN_548;
  wire  GEN_549;
  wire  GEN_550;
  wire  GEN_551;
  wire  GEN_552;
  wire  GEN_553;
  wire  GEN_554;
  wire  GEN_555;
  wire  GEN_556;
  wire  GEN_557;
  wire  GEN_558;
  wire  GEN_559;
  wire  GEN_560;
  wire  GEN_561;
  wire  GEN_562;
  wire  GEN_563;
  wire  GEN_564;
  wire  GEN_565;
  wire  GEN_566;
  wire  GEN_567;
  wire  GEN_568;
  wire  GEN_569;
  wire  GEN_570;
  wire  GEN_571;
  wire  GEN_572;
  wire  GEN_573;
  wire  GEN_574;
  wire  GEN_575;
  wire  GEN_576;
  wire  GEN_577;
  wire  GEN_578;
  wire  GEN_579;
  wire  GEN_580;
  wire  GEN_581;
  wire  GEN_582;
  wire  GEN_583;
  wire  GEN_584;
  wire  GEN_585;
  wire  GEN_586;
  wire  GEN_587;
  wire  GEN_588;
  wire  GEN_589;
  wire  GEN_590;
  wire  GEN_591;
  wire  GEN_592;
  wire  GEN_593;
  wire  GEN_594;
  wire  GEN_595;
  wire  GEN_596;
  wire  GEN_597;
  wire  GEN_598;
  wire  GEN_599;
  wire  GEN_600;
  wire  GEN_601;
  wire  GEN_602;
  wire  GEN_603;
  wire  GEN_604;
  wire  GEN_605;
  wire  GEN_606;
  wire  GEN_607;
  wire  GEN_608;
  wire  GEN_609;
  wire  GEN_610;
  wire  GEN_611;
  wire  GEN_612;
  wire  GEN_613;
  wire  GEN_614;
  wire  GEN_615;
  wire  GEN_616;
  wire  GEN_617;
  wire  GEN_618;
  wire  GEN_619;
  wire  GEN_620;
  wire  GEN_621;
  wire  GEN_622;
  wire  GEN_623;
  wire  GEN_624;
  wire  GEN_625;
  wire  GEN_626;
  wire  GEN_627;
  wire  GEN_628;
  wire  GEN_629;
  wire  GEN_630;
  wire  GEN_631;
  wire  GEN_632;
  wire  GEN_633;
  wire  GEN_634;
  wire  GEN_635;
  wire  GEN_636;
  wire  GEN_637;
  wire  GEN_638;
  wire  GEN_639;
  wire  GEN_640;
  wire  GEN_641;
  wire  GEN_642;
  wire  GEN_643;
  wire  GEN_644;
  wire  GEN_645;
  wire  GEN_646;
  wire  GEN_647;
  wire  GEN_648;
  wire  GEN_649;
  wire  GEN_650;
  wire  GEN_651;
  wire  GEN_652;
  wire  GEN_653;
  wire  GEN_654;
  wire  GEN_655;
  wire  GEN_656;
  wire  GEN_657;
  wire  GEN_658;
  wire  GEN_659;
  wire  GEN_660;
  wire  GEN_661;
  wire  GEN_662;
  wire  GEN_663;
  wire  GEN_664;
  wire  GEN_665;
  wire  GEN_666;
  wire  GEN_667;
  wire  GEN_668;
  wire  GEN_669;
  wire  GEN_670;
  wire  GEN_671;
  wire  GEN_672;
  wire  GEN_673;
  wire  GEN_674;
  wire  GEN_675;
  wire  GEN_676;
  wire  GEN_677;
  wire  GEN_678;
  wire  GEN_679;
  wire  GEN_680;
  wire  GEN_681;
  wire  GEN_682;
  wire  GEN_683;
  wire  GEN_684;
  wire  GEN_685;
  wire  GEN_686;
  wire  GEN_687;
  wire  GEN_688;
  wire  GEN_689;
  wire  GEN_690;
  wire  GEN_691;
  wire  GEN_692;
  wire  GEN_693;
  wire  GEN_694;
  wire  GEN_695;
  wire  GEN_696;
  wire  GEN_697;
  wire  GEN_698;
  wire  GEN_699;
  wire  GEN_700;
  wire  GEN_701;
  wire  GEN_702;
  wire  GEN_703;
  wire  GEN_704;
  wire  GEN_705;
  wire  GEN_706;
  wire  GEN_707;
  wire  GEN_708;
  wire  GEN_709;
  wire  GEN_710;
  wire  GEN_711;
  wire  GEN_712;
  wire  GEN_713;
  wire  GEN_714;
  wire  GEN_715;
  wire  GEN_716;
  wire  GEN_717;
  wire  GEN_718;
  wire  GEN_719;
  wire  GEN_720;
  wire  GEN_721;
  wire  GEN_722;
  wire  GEN_723;
  wire  GEN_724;
  wire  GEN_725;
  wire  GEN_726;
  wire  GEN_727;
  wire  GEN_728;
  wire  GEN_729;
  wire  GEN_730;
  wire  GEN_731;
  wire  GEN_732;
  wire  GEN_733;
  wire  GEN_734;
  wire  GEN_735;
  wire  GEN_736;
  wire  GEN_737;
  wire  GEN_738;
  wire  GEN_739;
  wire  GEN_740;
  wire  GEN_741;
  wire  GEN_742;
  wire  GEN_743;
  wire  GEN_744;
  wire  GEN_745;
  wire  GEN_746;
  wire  GEN_747;
  wire  GEN_748;
  wire  GEN_749;
  wire  GEN_750;
  wire  GEN_751;
  wire  GEN_752;
  wire  GEN_753;
  wire  GEN_754;
  wire  GEN_755;
  wire  GEN_756;
  wire  GEN_757;
  wire  GEN_758;
  wire  GEN_759;
  wire  GEN_760;
  wire  GEN_761;
  wire  GEN_762;
  wire  GEN_763;
  wire  GEN_764;
  wire  GEN_765;
  wire  GEN_766;
  wire  GEN_767;
  wire  GEN_768;
  wire  GEN_769;
  wire  GEN_770;
  wire  GEN_771;
  wire  GEN_772;
  wire  GEN_773;
  wire  GEN_774;
  wire  GEN_775;
  wire  GEN_776;
  wire  GEN_777;
  wire  GEN_778;
  wire  GEN_779;
  wire  GEN_780;
  wire  GEN_781;
  wire  GEN_782;
  wire  GEN_783;
  wire  GEN_784;
  wire  GEN_785;
  wire  GEN_786;
  wire  GEN_787;
  wire  GEN_788;
  wire  GEN_789;
  wire  GEN_790;
  wire  GEN_791;
  wire  GEN_792;
  wire  GEN_793;
  wire  GEN_794;
  wire  GEN_795;
  wire  GEN_796;
  wire  GEN_797;
  wire  GEN_798;
  wire  GEN_799;
  wire  GEN_800;
  wire  GEN_801;
  wire  GEN_802;
  wire  GEN_803;
  wire  GEN_804;
  wire  GEN_805;
  wire  GEN_806;
  wire  GEN_807;
  wire  GEN_808;
  wire  GEN_809;
  wire  GEN_810;
  wire  GEN_811;
  wire  GEN_812;
  wire  GEN_813;
  wire  GEN_814;
  wire  GEN_815;
  wire  GEN_816;
  wire  GEN_817;
  wire  GEN_818;
  wire  GEN_819;
  wire  GEN_820;
  wire  GEN_821;
  wire  GEN_822;
  wire  GEN_823;
  wire  GEN_824;
  wire  GEN_825;
  wire  GEN_826;
  wire  GEN_827;
  wire  GEN_828;
  wire  GEN_829;
  wire  GEN_830;
  wire  GEN_831;
  wire  GEN_832;
  wire  GEN_833;
  wire  GEN_834;
  wire  GEN_835;
  wire  GEN_836;
  wire  GEN_837;
  wire  GEN_838;
  wire  GEN_839;
  wire  GEN_840;
  wire  GEN_841;
  wire  GEN_842;
  wire  GEN_843;
  wire  GEN_844;
  wire  GEN_845;
  wire  GEN_846;
  wire  GEN_847;
  wire  GEN_848;
  wire  GEN_849;
  wire  GEN_850;
  wire  GEN_851;
  wire  GEN_852;
  wire  GEN_853;
  wire  GEN_854;
  wire  GEN_855;
  wire  GEN_856;
  wire  GEN_857;
  wire  GEN_858;
  wire  GEN_859;
  wire  GEN_860;
  wire  GEN_861;
  wire  GEN_862;
  wire  GEN_863;
  wire  GEN_864;
  wire  GEN_865;
  wire  GEN_866;
  wire  GEN_867;
  wire  GEN_868;
  wire  GEN_869;
  wire  GEN_870;
  wire  GEN_871;
  wire  GEN_872;
  wire  GEN_873;
  wire  GEN_874;
  wire  GEN_875;
  wire  GEN_876;
  wire  GEN_877;
  wire  GEN_878;
  wire  GEN_879;
  wire  GEN_880;
  wire  GEN_881;
  wire  GEN_882;
  wire  GEN_883;
  wire  GEN_884;
  wire  GEN_885;
  wire  GEN_886;
  wire  GEN_887;
  wire  GEN_888;
  wire  GEN_889;
  wire  GEN_890;
  wire  GEN_891;
  wire  GEN_892;
  wire  GEN_893;
  wire  GEN_894;
  wire  GEN_895;
  wire  GEN_896;
  wire  GEN_897;
  wire  GEN_898;
  wire  GEN_899;
  wire  GEN_900;
  wire  GEN_901;
  wire  GEN_902;
  wire  GEN_903;
  wire  GEN_904;
  wire  GEN_905;
  wire  GEN_906;
  wire  GEN_907;
  wire  GEN_908;
  wire  GEN_909;
  wire  GEN_910;
  wire  GEN_911;
  wire  GEN_912;
  wire  GEN_913;
  wire  GEN_914;
  wire  GEN_915;
  wire  GEN_916;
  wire  GEN_917;
  wire  GEN_918;
  wire  GEN_919;
  wire  GEN_920;
  wire  GEN_921;
  wire  GEN_922;
  wire  GEN_923;
  wire  GEN_924;
  wire  GEN_925;
  wire  GEN_926;
  wire  GEN_927;
  wire  GEN_928;
  wire  GEN_929;
  wire  GEN_930;
  wire  GEN_931;
  wire  GEN_932;
  wire  GEN_933;
  wire  GEN_4;
  wire  GEN_934;
  wire  GEN_935;
  wire  GEN_936;
  wire  GEN_937;
  wire  GEN_938;
  wire  GEN_939;
  wire  GEN_940;
  wire  GEN_941;
  wire  GEN_942;
  wire  GEN_943;
  wire  GEN_944;
  wire  GEN_945;
  wire  GEN_946;
  wire  GEN_947;
  wire  GEN_948;
  wire  GEN_949;
  wire  GEN_950;
  wire  GEN_951;
  wire  GEN_952;
  wire  GEN_953;
  wire  GEN_954;
  wire  GEN_955;
  wire  GEN_956;
  wire  GEN_957;
  wire  GEN_958;
  wire  GEN_959;
  wire  GEN_960;
  wire  GEN_961;
  wire  GEN_962;
  wire  GEN_963;
  wire  GEN_964;
  wire  GEN_965;
  wire  GEN_966;
  wire  GEN_967;
  wire  GEN_968;
  wire  GEN_969;
  wire  GEN_970;
  wire  GEN_971;
  wire  GEN_972;
  wire  GEN_973;
  wire  GEN_974;
  wire  GEN_975;
  wire  GEN_976;
  wire  GEN_977;
  wire  GEN_978;
  wire  GEN_979;
  wire  GEN_980;
  wire  GEN_981;
  wire  GEN_982;
  wire  GEN_983;
  wire  GEN_984;
  wire  GEN_985;
  wire  GEN_986;
  wire  GEN_987;
  wire  GEN_988;
  wire  GEN_989;
  wire  GEN_990;
  wire  GEN_991;
  wire  GEN_992;
  wire  GEN_993;
  wire  GEN_994;
  wire  GEN_995;
  wire  GEN_996;
  wire  GEN_997;
  wire  GEN_998;
  wire  GEN_999;
  wire  GEN_1000;
  wire  GEN_1001;
  wire  GEN_1002;
  wire  GEN_1003;
  wire  GEN_1004;
  wire  GEN_1005;
  wire  GEN_1006;
  wire  GEN_1007;
  wire  GEN_1008;
  wire  GEN_1009;
  wire  GEN_1010;
  wire  GEN_1011;
  wire  GEN_1012;
  wire  GEN_1013;
  wire  GEN_1014;
  wire  GEN_1015;
  wire  GEN_1016;
  wire  GEN_1017;
  wire  GEN_1018;
  wire  GEN_1019;
  wire  GEN_1020;
  wire  GEN_1021;
  wire  GEN_1022;
  wire  GEN_1023;
  wire  GEN_1024;
  wire  GEN_1025;
  wire  GEN_1026;
  wire  GEN_1027;
  wire  GEN_1028;
  wire  GEN_1029;
  wire  GEN_1030;
  wire  GEN_1031;
  wire  GEN_1032;
  wire  GEN_1033;
  wire  GEN_1034;
  wire  GEN_1035;
  wire  GEN_1036;
  wire  GEN_1037;
  wire  GEN_1038;
  wire  GEN_1039;
  wire  GEN_1040;
  wire  GEN_1041;
  wire  GEN_1042;
  wire  GEN_1043;
  wire  GEN_1044;
  wire  GEN_1045;
  wire  GEN_1046;
  wire  GEN_1047;
  wire  GEN_1048;
  wire  GEN_1049;
  wire  GEN_1050;
  wire  GEN_1051;
  wire  GEN_1052;
  wire  GEN_1053;
  wire  GEN_1054;
  wire  GEN_1055;
  wire  GEN_1056;
  wire  GEN_1057;
  wire  GEN_1058;
  wire  GEN_1059;
  wire  GEN_1060;
  wire  GEN_1061;
  wire  GEN_1062;
  wire  GEN_1063;
  wire  GEN_1064;
  wire  GEN_1065;
  wire  GEN_1066;
  wire  GEN_1067;
  wire  GEN_1068;
  wire  GEN_1069;
  wire  GEN_1070;
  wire  GEN_1071;
  wire  GEN_1072;
  wire  GEN_1073;
  wire  GEN_1074;
  wire  GEN_1075;
  wire  GEN_1076;
  wire  GEN_1077;
  wire  GEN_1078;
  wire  GEN_1079;
  wire  GEN_1080;
  wire  GEN_1081;
  wire  GEN_1082;
  wire  GEN_1083;
  wire  GEN_1084;
  wire  GEN_1085;
  wire  GEN_1086;
  wire  GEN_1087;
  wire  GEN_1088;
  wire  GEN_1089;
  wire  GEN_1090;
  wire  GEN_1091;
  wire  GEN_1092;
  wire  GEN_1093;
  wire  GEN_1094;
  wire  GEN_1095;
  wire  GEN_1096;
  wire  GEN_1097;
  wire  GEN_1098;
  wire  GEN_1099;
  wire  GEN_1100;
  wire  GEN_1101;
  wire  GEN_1102;
  wire  GEN_1103;
  wire  GEN_1104;
  wire  GEN_1105;
  wire  GEN_1106;
  wire  GEN_1107;
  wire  GEN_1108;
  wire  GEN_1109;
  wire  GEN_1110;
  wire  GEN_1111;
  wire  GEN_1112;
  wire  GEN_1113;
  wire  GEN_1114;
  wire  GEN_1115;
  wire  GEN_1116;
  wire  GEN_1117;
  wire  GEN_1118;
  wire  GEN_1119;
  wire  GEN_1120;
  wire  GEN_1121;
  wire  GEN_1122;
  wire  GEN_1123;
  wire  GEN_1124;
  wire  GEN_1125;
  wire  GEN_1126;
  wire  GEN_1127;
  wire  GEN_1128;
  wire  GEN_1129;
  wire  GEN_1130;
  wire  GEN_1131;
  wire  GEN_1132;
  wire  GEN_1133;
  wire  GEN_1134;
  wire  GEN_1135;
  wire  GEN_1136;
  wire  GEN_1137;
  wire  GEN_1138;
  wire  GEN_1139;
  wire  GEN_1140;
  wire  GEN_1141;
  wire  GEN_1142;
  wire  GEN_1143;
  wire  GEN_1144;
  wire  GEN_1145;
  wire  GEN_1146;
  wire  GEN_1147;
  wire  GEN_1148;
  wire  GEN_1149;
  wire  GEN_1150;
  wire  GEN_1151;
  wire  GEN_1152;
  wire  GEN_1153;
  wire  GEN_1154;
  wire  GEN_1155;
  wire  GEN_1156;
  wire  GEN_1157;
  wire  GEN_1158;
  wire  GEN_1159;
  wire  GEN_1160;
  wire  GEN_1161;
  wire  GEN_1162;
  wire  GEN_1163;
  wire  GEN_1164;
  wire  GEN_1165;
  wire  GEN_1166;
  wire  GEN_1167;
  wire  GEN_1168;
  wire  GEN_1169;
  wire  GEN_1170;
  wire  GEN_1171;
  wire  GEN_1172;
  wire  GEN_1173;
  wire  GEN_1174;
  wire  GEN_1175;
  wire  GEN_1176;
  wire  GEN_1177;
  wire  GEN_1178;
  wire  GEN_1179;
  wire  GEN_1180;
  wire  GEN_1181;
  wire  GEN_1182;
  wire  GEN_1183;
  wire  GEN_1184;
  wire  GEN_1185;
  wire  GEN_1186;
  wire  GEN_1187;
  wire  GEN_1188;
  wire  GEN_1189;
  wire  GEN_1190;
  wire  GEN_1191;
  wire  GEN_1192;
  wire  GEN_1193;
  wire  GEN_1194;
  wire  GEN_1195;
  wire  GEN_1196;
  wire  GEN_1197;
  wire  GEN_1198;
  wire  GEN_1199;
  wire  GEN_1200;
  wire  GEN_1201;
  wire  GEN_1202;
  wire  GEN_1203;
  wire  GEN_1204;
  wire  GEN_1205;
  wire  GEN_1206;
  wire  GEN_1207;
  wire  GEN_1208;
  wire  GEN_1209;
  wire  GEN_1210;
  wire  GEN_1211;
  wire  GEN_1212;
  wire  GEN_1213;
  wire  GEN_1214;
  wire  GEN_1215;
  wire  GEN_1216;
  wire  GEN_1217;
  wire  GEN_1218;
  wire  GEN_1219;
  wire  GEN_1220;
  wire  GEN_1221;
  wire  GEN_1222;
  wire  GEN_1223;
  wire  GEN_1224;
  wire  GEN_1225;
  wire  GEN_1226;
  wire  GEN_1227;
  wire  GEN_1228;
  wire  GEN_1229;
  wire  GEN_1230;
  wire  GEN_1231;
  wire  GEN_1232;
  wire  GEN_1233;
  wire  GEN_1234;
  wire  GEN_1235;
  wire  GEN_1236;
  wire  GEN_1237;
  wire  GEN_1238;
  wire  GEN_1239;
  wire  GEN_1240;
  wire  GEN_1241;
  wire  GEN_1242;
  wire  GEN_1243;
  wire  GEN_1244;
  wire  GEN_1245;
  wire  GEN_1246;
  wire  GEN_1247;
  wire  GEN_1248;
  wire  GEN_1249;
  wire  GEN_1250;
  wire  GEN_1251;
  wire  GEN_1252;
  wire  GEN_1253;
  wire  GEN_1254;
  wire  GEN_1255;
  wire  GEN_1256;
  wire  GEN_1257;
  wire  GEN_1258;
  wire  GEN_1259;
  wire  GEN_1260;
  wire  GEN_1261;
  wire  GEN_1262;
  wire  GEN_1263;
  wire  GEN_1264;
  wire  GEN_1265;
  wire  GEN_1266;
  wire  GEN_1267;
  wire  GEN_1268;
  wire  GEN_1269;
  wire  GEN_1270;
  wire  GEN_1271;
  wire  GEN_1272;
  wire  GEN_1273;
  wire  GEN_1274;
  wire  GEN_1275;
  wire  GEN_1276;
  wire  GEN_1277;
  wire  GEN_1278;
  wire  GEN_1279;
  wire  GEN_1280;
  wire  GEN_1281;
  wire  GEN_1282;
  wire  GEN_1283;
  wire  GEN_1284;
  wire  GEN_1285;
  wire  GEN_1286;
  wire  GEN_1287;
  wire  GEN_1288;
  wire  GEN_1289;
  wire  GEN_1290;
  wire  GEN_1291;
  wire  GEN_1292;
  wire  GEN_1293;
  wire  GEN_1294;
  wire  GEN_1295;
  wire  GEN_1296;
  wire  GEN_1297;
  wire  GEN_1298;
  wire  GEN_1299;
  wire  GEN_1300;
  wire  GEN_1301;
  wire  GEN_1302;
  wire  GEN_1303;
  wire  GEN_1304;
  wire  GEN_1305;
  wire  GEN_1306;
  wire  GEN_1307;
  wire  GEN_1308;
  wire  GEN_1309;
  wire  GEN_1310;
  wire  GEN_1311;
  wire  GEN_1312;
  wire  GEN_1313;
  wire  GEN_1314;
  wire  GEN_1315;
  wire  GEN_1316;
  wire  GEN_1317;
  wire  GEN_1318;
  wire  GEN_1319;
  wire  GEN_1320;
  wire  GEN_1321;
  wire  GEN_1322;
  wire  GEN_1323;
  wire  GEN_1324;
  wire  GEN_1325;
  wire  GEN_1326;
  wire  GEN_1327;
  wire  GEN_1328;
  wire  GEN_1329;
  wire  GEN_1330;
  wire  GEN_1331;
  wire  GEN_1332;
  wire  GEN_1333;
  wire  GEN_1334;
  wire  GEN_1335;
  wire  GEN_1336;
  wire  GEN_1337;
  wire  GEN_1338;
  wire  GEN_1339;
  wire  GEN_1340;
  wire  GEN_1341;
  wire  GEN_1342;
  wire  GEN_1343;
  wire  GEN_1344;
  wire  GEN_1345;
  wire  GEN_1346;
  wire  GEN_1347;
  wire  GEN_1348;
  wire  GEN_1349;
  wire  GEN_1350;
  wire  GEN_1351;
  wire  GEN_1352;
  wire  GEN_1353;
  wire  GEN_1354;
  wire  GEN_1355;
  wire  GEN_1356;
  wire  GEN_1357;
  wire  GEN_1358;
  wire  GEN_1359;
  wire  GEN_1360;
  wire  GEN_1361;
  wire  GEN_1362;
  wire  GEN_1363;
  wire  GEN_1364;
  wire  GEN_1365;
  wire  GEN_1366;
  wire  GEN_1367;
  wire  GEN_1368;
  wire  GEN_1369;
  wire  GEN_1370;
  wire  GEN_1371;
  wire  GEN_1372;
  wire  GEN_1373;
  wire  GEN_1374;
  wire  GEN_1375;
  wire  GEN_1376;
  wire  GEN_1377;
  wire  GEN_1378;
  wire  GEN_1379;
  wire  GEN_1380;
  wire  GEN_1381;
  wire  GEN_1382;
  wire  GEN_1383;
  wire  GEN_1384;
  wire  GEN_1385;
  wire  GEN_1386;
  wire  GEN_1387;
  wire  GEN_1388;
  wire  GEN_1389;
  wire  GEN_1390;
  wire  GEN_1391;
  wire  GEN_1392;
  wire  GEN_1393;
  wire  GEN_1394;
  wire  GEN_1395;
  wire  GEN_1396;
  wire  GEN_1397;
  wire  GEN_1398;
  wire  GEN_1399;
  wire  GEN_1400;
  wire  GEN_1401;
  wire  GEN_1402;
  wire  GEN_1403;
  wire  GEN_1404;
  wire  GEN_1405;
  wire  GEN_1406;
  wire  GEN_1407;
  wire  GEN_1408;
  wire  GEN_1409;
  wire  GEN_1410;
  wire  GEN_1411;
  wire  GEN_1412;
  wire  GEN_1413;
  wire  GEN_1414;
  wire  GEN_1415;
  wire  GEN_1416;
  wire  GEN_1417;
  wire  GEN_1418;
  wire  GEN_1419;
  wire  GEN_1420;
  wire  GEN_1421;
  wire  GEN_1422;
  wire  GEN_1423;
  wire  GEN_1424;
  wire  GEN_1425;
  wire  GEN_1426;
  wire  GEN_1427;
  wire  GEN_1428;
  wire  GEN_1429;
  wire  GEN_1430;
  wire  GEN_1431;
  wire  GEN_1432;
  wire  GEN_1433;
  wire  GEN_1434;
  wire  GEN_1435;
  wire  GEN_1436;
  wire  GEN_1437;
  wire  GEN_1438;
  wire  GEN_1439;
  wire  GEN_1440;
  wire  GEN_1441;
  wire  GEN_1442;
  wire  GEN_1443;
  wire  GEN_1444;
  wire  T_24257;
  wire  GEN_5;
  wire  GEN_1445;
  wire  GEN_1446;
  wire  GEN_1447;
  wire  GEN_1448;
  wire  GEN_1449;
  wire  GEN_1450;
  wire  GEN_1451;
  wire  GEN_1452;
  wire  GEN_1453;
  wire  GEN_1454;
  wire  GEN_1455;
  wire  GEN_1456;
  wire  GEN_1457;
  wire  GEN_1458;
  wire  GEN_1459;
  wire  GEN_1460;
  wire  GEN_1461;
  wire  GEN_1462;
  wire  GEN_1463;
  wire  GEN_1464;
  wire  GEN_1465;
  wire  GEN_1466;
  wire  GEN_1467;
  wire  GEN_1468;
  wire  GEN_1469;
  wire  GEN_1470;
  wire  GEN_1471;
  wire  GEN_1472;
  wire  GEN_1473;
  wire  GEN_1474;
  wire  GEN_1475;
  wire  GEN_1476;
  wire  GEN_1477;
  wire  GEN_1478;
  wire  GEN_1479;
  wire  GEN_1480;
  wire  GEN_1481;
  wire  GEN_1482;
  wire  GEN_1483;
  wire  GEN_1484;
  wire  GEN_1485;
  wire  GEN_1486;
  wire  GEN_1487;
  wire  GEN_1488;
  wire  GEN_1489;
  wire  GEN_1490;
  wire  GEN_1491;
  wire  GEN_1492;
  wire  GEN_1493;
  wire  GEN_1494;
  wire  GEN_1495;
  wire  GEN_1496;
  wire  GEN_1497;
  wire  GEN_1498;
  wire  GEN_1499;
  wire  GEN_1500;
  wire  GEN_1501;
  wire  GEN_1502;
  wire  GEN_1503;
  wire  GEN_1504;
  wire  GEN_1505;
  wire  GEN_1506;
  wire  GEN_1507;
  wire  GEN_1508;
  wire  GEN_1509;
  wire  GEN_1510;
  wire  GEN_1511;
  wire  GEN_1512;
  wire  GEN_1513;
  wire  GEN_1514;
  wire  GEN_1515;
  wire  GEN_1516;
  wire  GEN_1517;
  wire  GEN_1518;
  wire  GEN_1519;
  wire  GEN_1520;
  wire  GEN_1521;
  wire  GEN_1522;
  wire  GEN_1523;
  wire  GEN_1524;
  wire  GEN_1525;
  wire  GEN_1526;
  wire  GEN_1527;
  wire  GEN_1528;
  wire  GEN_1529;
  wire  GEN_1530;
  wire  GEN_1531;
  wire  GEN_1532;
  wire  GEN_1533;
  wire  GEN_1534;
  wire  GEN_1535;
  wire  GEN_1536;
  wire  GEN_1537;
  wire  GEN_1538;
  wire  GEN_1539;
  wire  GEN_1540;
  wire  GEN_1541;
  wire  GEN_1542;
  wire  GEN_1543;
  wire  GEN_1544;
  wire  GEN_1545;
  wire  GEN_1546;
  wire  GEN_1547;
  wire  GEN_1548;
  wire  GEN_1549;
  wire  GEN_1550;
  wire  GEN_1551;
  wire  GEN_1552;
  wire  GEN_1553;
  wire  GEN_1554;
  wire  GEN_1555;
  wire  GEN_1556;
  wire  GEN_1557;
  wire  GEN_1558;
  wire  GEN_1559;
  wire  GEN_1560;
  wire  GEN_1561;
  wire  GEN_1562;
  wire  GEN_1563;
  wire  GEN_1564;
  wire  GEN_1565;
  wire  GEN_1566;
  wire  GEN_1567;
  wire  GEN_1568;
  wire  GEN_1569;
  wire  GEN_1570;
  wire  GEN_1571;
  wire  GEN_1572;
  wire  GEN_1573;
  wire  GEN_1574;
  wire  GEN_1575;
  wire  GEN_1576;
  wire  GEN_1577;
  wire  GEN_1578;
  wire  GEN_1579;
  wire  GEN_1580;
  wire  GEN_1581;
  wire  GEN_1582;
  wire  GEN_1583;
  wire  GEN_1584;
  wire  GEN_1585;
  wire  GEN_1586;
  wire  GEN_1587;
  wire  GEN_1588;
  wire  GEN_1589;
  wire  GEN_1590;
  wire  GEN_1591;
  wire  GEN_1592;
  wire  GEN_1593;
  wire  GEN_1594;
  wire  GEN_1595;
  wire  GEN_1596;
  wire  GEN_1597;
  wire  GEN_1598;
  wire  GEN_1599;
  wire  GEN_1600;
  wire  GEN_1601;
  wire  GEN_1602;
  wire  GEN_1603;
  wire  GEN_1604;
  wire  GEN_1605;
  wire  GEN_1606;
  wire  GEN_1607;
  wire  GEN_1608;
  wire  GEN_1609;
  wire  GEN_1610;
  wire  GEN_1611;
  wire  GEN_1612;
  wire  GEN_1613;
  wire  GEN_1614;
  wire  GEN_1615;
  wire  GEN_1616;
  wire  GEN_1617;
  wire  GEN_1618;
  wire  GEN_1619;
  wire  GEN_1620;
  wire  GEN_1621;
  wire  GEN_1622;
  wire  GEN_1623;
  wire  GEN_1624;
  wire  GEN_1625;
  wire  GEN_1626;
  wire  GEN_1627;
  wire  GEN_1628;
  wire  GEN_1629;
  wire  GEN_1630;
  wire  GEN_1631;
  wire  GEN_1632;
  wire  GEN_1633;
  wire  GEN_1634;
  wire  GEN_1635;
  wire  GEN_1636;
  wire  GEN_1637;
  wire  GEN_1638;
  wire  GEN_1639;
  wire  GEN_1640;
  wire  GEN_1641;
  wire  GEN_1642;
  wire  GEN_1643;
  wire  GEN_1644;
  wire  GEN_1645;
  wire  GEN_1646;
  wire  GEN_1647;
  wire  GEN_1648;
  wire  GEN_1649;
  wire  GEN_1650;
  wire  GEN_1651;
  wire  GEN_1652;
  wire  GEN_1653;
  wire  GEN_1654;
  wire  GEN_1655;
  wire  GEN_1656;
  wire  GEN_1657;
  wire  GEN_1658;
  wire  GEN_1659;
  wire  GEN_1660;
  wire  GEN_1661;
  wire  GEN_1662;
  wire  GEN_1663;
  wire  GEN_1664;
  wire  GEN_1665;
  wire  GEN_1666;
  wire  GEN_1667;
  wire  GEN_1668;
  wire  GEN_1669;
  wire  GEN_1670;
  wire  GEN_1671;
  wire  GEN_1672;
  wire  GEN_1673;
  wire  GEN_1674;
  wire  GEN_1675;
  wire  GEN_1676;
  wire  GEN_1677;
  wire  GEN_1678;
  wire  GEN_1679;
  wire  GEN_1680;
  wire  GEN_1681;
  wire  GEN_1682;
  wire  GEN_1683;
  wire  GEN_1684;
  wire  GEN_1685;
  wire  GEN_1686;
  wire  GEN_1687;
  wire  GEN_1688;
  wire  GEN_1689;
  wire  GEN_1690;
  wire  GEN_1691;
  wire  GEN_1692;
  wire  GEN_1693;
  wire  GEN_1694;
  wire  GEN_1695;
  wire  GEN_1696;
  wire  GEN_1697;
  wire  GEN_1698;
  wire  GEN_1699;
  wire  GEN_1700;
  wire  GEN_1701;
  wire  GEN_1702;
  wire  GEN_1703;
  wire  GEN_1704;
  wire  GEN_1705;
  wire  GEN_1706;
  wire  GEN_1707;
  wire  GEN_1708;
  wire  GEN_1709;
  wire  GEN_1710;
  wire  GEN_1711;
  wire  GEN_1712;
  wire  GEN_1713;
  wire  GEN_1714;
  wire  GEN_1715;
  wire  GEN_1716;
  wire  GEN_1717;
  wire  GEN_1718;
  wire  GEN_1719;
  wire  GEN_1720;
  wire  GEN_1721;
  wire  GEN_1722;
  wire  GEN_1723;
  wire  GEN_1724;
  wire  GEN_1725;
  wire  GEN_1726;
  wire  GEN_1727;
  wire  GEN_1728;
  wire  GEN_1729;
  wire  GEN_1730;
  wire  GEN_1731;
  wire  GEN_1732;
  wire  GEN_1733;
  wire  GEN_1734;
  wire  GEN_1735;
  wire  GEN_1736;
  wire  GEN_1737;
  wire  GEN_1738;
  wire  GEN_1739;
  wire  GEN_1740;
  wire  GEN_1741;
  wire  GEN_1742;
  wire  GEN_1743;
  wire  GEN_1744;
  wire  GEN_1745;
  wire  GEN_1746;
  wire  GEN_1747;
  wire  GEN_1748;
  wire  GEN_1749;
  wire  GEN_1750;
  wire  GEN_1751;
  wire  GEN_1752;
  wire  GEN_1753;
  wire  GEN_1754;
  wire  GEN_1755;
  wire  GEN_1756;
  wire  GEN_1757;
  wire  GEN_1758;
  wire  GEN_1759;
  wire  GEN_1760;
  wire  GEN_1761;
  wire  GEN_1762;
  wire  GEN_1763;
  wire  GEN_1764;
  wire  GEN_1765;
  wire  GEN_1766;
  wire  GEN_1767;
  wire  GEN_1768;
  wire  GEN_1769;
  wire  GEN_1770;
  wire  GEN_1771;
  wire  GEN_1772;
  wire  GEN_1773;
  wire  GEN_1774;
  wire  GEN_1775;
  wire  GEN_1776;
  wire  GEN_1777;
  wire  GEN_1778;
  wire  GEN_1779;
  wire  GEN_1780;
  wire  GEN_1781;
  wire  GEN_1782;
  wire  GEN_1783;
  wire  GEN_1784;
  wire  GEN_1785;
  wire  GEN_1786;
  wire  GEN_1787;
  wire  GEN_1788;
  wire  GEN_1789;
  wire  GEN_1790;
  wire  GEN_1791;
  wire  GEN_1792;
  wire  GEN_1793;
  wire  GEN_1794;
  wire  GEN_1795;
  wire  GEN_1796;
  wire  GEN_1797;
  wire  GEN_1798;
  wire  GEN_1799;
  wire  GEN_1800;
  wire  GEN_1801;
  wire  GEN_1802;
  wire  GEN_1803;
  wire  GEN_1804;
  wire  GEN_1805;
  wire  GEN_1806;
  wire  GEN_1807;
  wire  GEN_1808;
  wire  GEN_1809;
  wire  GEN_1810;
  wire  GEN_1811;
  wire  GEN_1812;
  wire  GEN_1813;
  wire  GEN_1814;
  wire  GEN_1815;
  wire  GEN_1816;
  wire  GEN_1817;
  wire  GEN_1818;
  wire  GEN_1819;
  wire  GEN_1820;
  wire  GEN_1821;
  wire  GEN_1822;
  wire  GEN_1823;
  wire  GEN_1824;
  wire  GEN_1825;
  wire  GEN_1826;
  wire  GEN_1827;
  wire  GEN_1828;
  wire  GEN_1829;
  wire  GEN_1830;
  wire  GEN_1831;
  wire  GEN_1832;
  wire  GEN_1833;
  wire  GEN_1834;
  wire  GEN_1835;
  wire  GEN_1836;
  wire  GEN_1837;
  wire  GEN_1838;
  wire  GEN_1839;
  wire  GEN_1840;
  wire  GEN_1841;
  wire  GEN_1842;
  wire  GEN_1843;
  wire  GEN_1844;
  wire  GEN_1845;
  wire  GEN_1846;
  wire  GEN_1847;
  wire  GEN_1848;
  wire  GEN_1849;
  wire  GEN_1850;
  wire  GEN_1851;
  wire  GEN_1852;
  wire  GEN_1853;
  wire  GEN_1854;
  wire  GEN_1855;
  wire  GEN_1856;
  wire  GEN_1857;
  wire  GEN_1858;
  wire  GEN_1859;
  wire  GEN_1860;
  wire  GEN_1861;
  wire  GEN_1862;
  wire  GEN_1863;
  wire  GEN_1864;
  wire  GEN_1865;
  wire  GEN_1866;
  wire  GEN_1867;
  wire  GEN_1868;
  wire  GEN_1869;
  wire  GEN_1870;
  wire  GEN_1871;
  wire  GEN_1872;
  wire  GEN_1873;
  wire  GEN_1874;
  wire  GEN_1875;
  wire  GEN_1876;
  wire  GEN_1877;
  wire  GEN_1878;
  wire  GEN_1879;
  wire  GEN_1880;
  wire  GEN_1881;
  wire  GEN_1882;
  wire  GEN_1883;
  wire  GEN_1884;
  wire  GEN_1885;
  wire  GEN_1886;
  wire  GEN_1887;
  wire  GEN_1888;
  wire  GEN_1889;
  wire  GEN_1890;
  wire  GEN_1891;
  wire  GEN_1892;
  wire  GEN_1893;
  wire  GEN_1894;
  wire  GEN_1895;
  wire  GEN_1896;
  wire  GEN_1897;
  wire  GEN_1898;
  wire  GEN_1899;
  wire  GEN_1900;
  wire  GEN_1901;
  wire  GEN_1902;
  wire  GEN_1903;
  wire  GEN_1904;
  wire  GEN_1905;
  wire  GEN_1906;
  wire  GEN_1907;
  wire  GEN_1908;
  wire  GEN_1909;
  wire  GEN_1910;
  wire  GEN_1911;
  wire  GEN_1912;
  wire  GEN_1913;
  wire  GEN_1914;
  wire  GEN_1915;
  wire  GEN_1916;
  wire  GEN_1917;
  wire  GEN_1918;
  wire  GEN_1919;
  wire  GEN_1920;
  wire  GEN_1921;
  wire  GEN_1922;
  wire  GEN_1923;
  wire  GEN_1924;
  wire  GEN_1925;
  wire  GEN_1926;
  wire  GEN_1927;
  wire  GEN_1928;
  wire  GEN_1929;
  wire  GEN_1930;
  wire  GEN_1931;
  wire  GEN_1932;
  wire  GEN_1933;
  wire  GEN_1934;
  wire  GEN_1935;
  wire  GEN_1936;
  wire  GEN_1937;
  wire  GEN_1938;
  wire  GEN_1939;
  wire  GEN_1940;
  wire  GEN_1941;
  wire  GEN_1942;
  wire  GEN_1943;
  wire  GEN_1944;
  wire  GEN_1945;
  wire  GEN_1946;
  wire  GEN_1947;
  wire  GEN_1948;
  wire  GEN_1949;
  wire  GEN_1950;
  wire  GEN_1951;
  wire  GEN_1952;
  wire  GEN_1953;
  wire  GEN_1954;
  wire  GEN_1955;
  wire  GEN_6;
  wire  GEN_1956;
  wire  GEN_1957;
  wire  GEN_1958;
  wire  GEN_1959;
  wire  GEN_1960;
  wire  GEN_1961;
  wire  GEN_1962;
  wire  GEN_1963;
  wire  GEN_1964;
  wire  GEN_1965;
  wire  GEN_1966;
  wire  GEN_1967;
  wire  GEN_1968;
  wire  GEN_1969;
  wire  GEN_1970;
  wire  GEN_1971;
  wire  GEN_1972;
  wire  GEN_1973;
  wire  GEN_1974;
  wire  GEN_1975;
  wire  GEN_1976;
  wire  GEN_1977;
  wire  GEN_1978;
  wire  GEN_1979;
  wire  GEN_1980;
  wire  GEN_1981;
  wire  GEN_1982;
  wire  GEN_1983;
  wire  GEN_1984;
  wire  GEN_1985;
  wire  GEN_1986;
  wire  GEN_1987;
  wire  GEN_1988;
  wire  GEN_1989;
  wire  GEN_1990;
  wire  GEN_1991;
  wire  GEN_1992;
  wire  GEN_1993;
  wire  GEN_1994;
  wire  GEN_1995;
  wire  GEN_1996;
  wire  GEN_1997;
  wire  GEN_1998;
  wire  GEN_1999;
  wire  GEN_2000;
  wire  GEN_2001;
  wire  GEN_2002;
  wire  GEN_2003;
  wire  GEN_2004;
  wire  GEN_2005;
  wire  GEN_2006;
  wire  GEN_2007;
  wire  GEN_2008;
  wire  GEN_2009;
  wire  GEN_2010;
  wire  GEN_2011;
  wire  GEN_2012;
  wire  GEN_2013;
  wire  GEN_2014;
  wire  GEN_2015;
  wire  GEN_2016;
  wire  GEN_2017;
  wire  GEN_2018;
  wire  GEN_2019;
  wire  GEN_2020;
  wire  GEN_2021;
  wire  GEN_2022;
  wire  GEN_2023;
  wire  GEN_2024;
  wire  GEN_2025;
  wire  GEN_2026;
  wire  GEN_2027;
  wire  GEN_2028;
  wire  GEN_2029;
  wire  GEN_2030;
  wire  GEN_2031;
  wire  GEN_2032;
  wire  GEN_2033;
  wire  GEN_2034;
  wire  GEN_2035;
  wire  GEN_2036;
  wire  GEN_2037;
  wire  GEN_2038;
  wire  GEN_2039;
  wire  GEN_2040;
  wire  GEN_2041;
  wire  GEN_2042;
  wire  GEN_2043;
  wire  GEN_2044;
  wire  GEN_2045;
  wire  GEN_2046;
  wire  GEN_2047;
  wire  GEN_2048;
  wire  GEN_2049;
  wire  GEN_2050;
  wire  GEN_2051;
  wire  GEN_2052;
  wire  GEN_2053;
  wire  GEN_2054;
  wire  GEN_2055;
  wire  GEN_2056;
  wire  GEN_2057;
  wire  GEN_2058;
  wire  GEN_2059;
  wire  GEN_2060;
  wire  GEN_2061;
  wire  GEN_2062;
  wire  GEN_2063;
  wire  GEN_2064;
  wire  GEN_2065;
  wire  GEN_2066;
  wire  GEN_2067;
  wire  GEN_2068;
  wire  GEN_2069;
  wire  GEN_2070;
  wire  GEN_2071;
  wire  GEN_2072;
  wire  GEN_2073;
  wire  GEN_2074;
  wire  GEN_2075;
  wire  GEN_2076;
  wire  GEN_2077;
  wire  GEN_2078;
  wire  GEN_2079;
  wire  GEN_2080;
  wire  GEN_2081;
  wire  GEN_2082;
  wire  GEN_2083;
  wire  GEN_2084;
  wire  GEN_2085;
  wire  GEN_2086;
  wire  GEN_2087;
  wire  GEN_2088;
  wire  GEN_2089;
  wire  GEN_2090;
  wire  GEN_2091;
  wire  GEN_2092;
  wire  GEN_2093;
  wire  GEN_2094;
  wire  GEN_2095;
  wire  GEN_2096;
  wire  GEN_2097;
  wire  GEN_2098;
  wire  GEN_2099;
  wire  GEN_2100;
  wire  GEN_2101;
  wire  GEN_2102;
  wire  GEN_2103;
  wire  GEN_2104;
  wire  GEN_2105;
  wire  GEN_2106;
  wire  GEN_2107;
  wire  GEN_2108;
  wire  GEN_2109;
  wire  GEN_2110;
  wire  GEN_2111;
  wire  GEN_2112;
  wire  GEN_2113;
  wire  GEN_2114;
  wire  GEN_2115;
  wire  GEN_2116;
  wire  GEN_2117;
  wire  GEN_2118;
  wire  GEN_2119;
  wire  GEN_2120;
  wire  GEN_2121;
  wire  GEN_2122;
  wire  GEN_2123;
  wire  GEN_2124;
  wire  GEN_2125;
  wire  GEN_2126;
  wire  GEN_2127;
  wire  GEN_2128;
  wire  GEN_2129;
  wire  GEN_2130;
  wire  GEN_2131;
  wire  GEN_2132;
  wire  GEN_2133;
  wire  GEN_2134;
  wire  GEN_2135;
  wire  GEN_2136;
  wire  GEN_2137;
  wire  GEN_2138;
  wire  GEN_2139;
  wire  GEN_2140;
  wire  GEN_2141;
  wire  GEN_2142;
  wire  GEN_2143;
  wire  GEN_2144;
  wire  GEN_2145;
  wire  GEN_2146;
  wire  GEN_2147;
  wire  GEN_2148;
  wire  GEN_2149;
  wire  GEN_2150;
  wire  GEN_2151;
  wire  GEN_2152;
  wire  GEN_2153;
  wire  GEN_2154;
  wire  GEN_2155;
  wire  GEN_2156;
  wire  GEN_2157;
  wire  GEN_2158;
  wire  GEN_2159;
  wire  GEN_2160;
  wire  GEN_2161;
  wire  GEN_2162;
  wire  GEN_2163;
  wire  GEN_2164;
  wire  GEN_2165;
  wire  GEN_2166;
  wire  GEN_2167;
  wire  GEN_2168;
  wire  GEN_2169;
  wire  GEN_2170;
  wire  GEN_2171;
  wire  GEN_2172;
  wire  GEN_2173;
  wire  GEN_2174;
  wire  GEN_2175;
  wire  GEN_2176;
  wire  GEN_2177;
  wire  GEN_2178;
  wire  GEN_2179;
  wire  GEN_2180;
  wire  GEN_2181;
  wire  GEN_2182;
  wire  GEN_2183;
  wire  GEN_2184;
  wire  GEN_2185;
  wire  GEN_2186;
  wire  GEN_2187;
  wire  GEN_2188;
  wire  GEN_2189;
  wire  GEN_2190;
  wire  GEN_2191;
  wire  GEN_2192;
  wire  GEN_2193;
  wire  GEN_2194;
  wire  GEN_2195;
  wire  GEN_2196;
  wire  GEN_2197;
  wire  GEN_2198;
  wire  GEN_2199;
  wire  GEN_2200;
  wire  GEN_2201;
  wire  GEN_2202;
  wire  GEN_2203;
  wire  GEN_2204;
  wire  GEN_2205;
  wire  GEN_2206;
  wire  GEN_2207;
  wire  GEN_2208;
  wire  GEN_2209;
  wire  GEN_2210;
  wire  GEN_2211;
  wire  GEN_2212;
  wire  GEN_2213;
  wire  GEN_2214;
  wire  GEN_2215;
  wire  GEN_2216;
  wire  GEN_2217;
  wire  GEN_2218;
  wire  GEN_2219;
  wire  GEN_2220;
  wire  GEN_2221;
  wire  GEN_2222;
  wire  GEN_2223;
  wire  GEN_2224;
  wire  GEN_2225;
  wire  GEN_2226;
  wire  GEN_2227;
  wire  GEN_2228;
  wire  GEN_2229;
  wire  GEN_2230;
  wire  GEN_2231;
  wire  GEN_2232;
  wire  GEN_2233;
  wire  GEN_2234;
  wire  GEN_2235;
  wire  GEN_2236;
  wire  GEN_2237;
  wire  GEN_2238;
  wire  GEN_2239;
  wire  GEN_2240;
  wire  GEN_2241;
  wire  GEN_2242;
  wire  GEN_2243;
  wire  GEN_2244;
  wire  GEN_2245;
  wire  GEN_2246;
  wire  GEN_2247;
  wire  GEN_2248;
  wire  GEN_2249;
  wire  GEN_2250;
  wire  GEN_2251;
  wire  GEN_2252;
  wire  GEN_2253;
  wire  GEN_2254;
  wire  GEN_2255;
  wire  GEN_2256;
  wire  GEN_2257;
  wire  GEN_2258;
  wire  GEN_2259;
  wire  GEN_2260;
  wire  GEN_2261;
  wire  GEN_2262;
  wire  GEN_2263;
  wire  GEN_2264;
  wire  GEN_2265;
  wire  GEN_2266;
  wire  GEN_2267;
  wire  GEN_2268;
  wire  GEN_2269;
  wire  GEN_2270;
  wire  GEN_2271;
  wire  GEN_2272;
  wire  GEN_2273;
  wire  GEN_2274;
  wire  GEN_2275;
  wire  GEN_2276;
  wire  GEN_2277;
  wire  GEN_2278;
  wire  GEN_2279;
  wire  GEN_2280;
  wire  GEN_2281;
  wire  GEN_2282;
  wire  GEN_2283;
  wire  GEN_2284;
  wire  GEN_2285;
  wire  GEN_2286;
  wire  GEN_2287;
  wire  GEN_2288;
  wire  GEN_2289;
  wire  GEN_2290;
  wire  GEN_2291;
  wire  GEN_2292;
  wire  GEN_2293;
  wire  GEN_2294;
  wire  GEN_2295;
  wire  GEN_2296;
  wire  GEN_2297;
  wire  GEN_2298;
  wire  GEN_2299;
  wire  GEN_2300;
  wire  GEN_2301;
  wire  GEN_2302;
  wire  GEN_2303;
  wire  GEN_2304;
  wire  GEN_2305;
  wire  GEN_2306;
  wire  GEN_2307;
  wire  GEN_2308;
  wire  GEN_2309;
  wire  GEN_2310;
  wire  GEN_2311;
  wire  GEN_2312;
  wire  GEN_2313;
  wire  GEN_2314;
  wire  GEN_2315;
  wire  GEN_2316;
  wire  GEN_2317;
  wire  GEN_2318;
  wire  GEN_2319;
  wire  GEN_2320;
  wire  GEN_2321;
  wire  GEN_2322;
  wire  GEN_2323;
  wire  GEN_2324;
  wire  GEN_2325;
  wire  GEN_2326;
  wire  GEN_2327;
  wire  GEN_2328;
  wire  GEN_2329;
  wire  GEN_2330;
  wire  GEN_2331;
  wire  GEN_2332;
  wire  GEN_2333;
  wire  GEN_2334;
  wire  GEN_2335;
  wire  GEN_2336;
  wire  GEN_2337;
  wire  GEN_2338;
  wire  GEN_2339;
  wire  GEN_2340;
  wire  GEN_2341;
  wire  GEN_2342;
  wire  GEN_2343;
  wire  GEN_2344;
  wire  GEN_2345;
  wire  GEN_2346;
  wire  GEN_2347;
  wire  GEN_2348;
  wire  GEN_2349;
  wire  GEN_2350;
  wire  GEN_2351;
  wire  GEN_2352;
  wire  GEN_2353;
  wire  GEN_2354;
  wire  GEN_2355;
  wire  GEN_2356;
  wire  GEN_2357;
  wire  GEN_2358;
  wire  GEN_2359;
  wire  GEN_2360;
  wire  GEN_2361;
  wire  GEN_2362;
  wire  GEN_2363;
  wire  GEN_2364;
  wire  GEN_2365;
  wire  GEN_2366;
  wire  GEN_2367;
  wire  GEN_2368;
  wire  GEN_2369;
  wire  GEN_2370;
  wire  GEN_2371;
  wire  GEN_2372;
  wire  GEN_2373;
  wire  GEN_2374;
  wire  GEN_2375;
  wire  GEN_2376;
  wire  GEN_2377;
  wire  GEN_2378;
  wire  GEN_2379;
  wire  GEN_2380;
  wire  GEN_2381;
  wire  GEN_2382;
  wire  GEN_2383;
  wire  GEN_2384;
  wire  GEN_2385;
  wire  GEN_2386;
  wire  GEN_2387;
  wire  GEN_2388;
  wire  GEN_2389;
  wire  GEN_2390;
  wire  GEN_2391;
  wire  GEN_2392;
  wire  GEN_2393;
  wire  GEN_2394;
  wire  GEN_2395;
  wire  GEN_2396;
  wire  GEN_2397;
  wire  GEN_2398;
  wire  GEN_2399;
  wire  GEN_2400;
  wire  GEN_2401;
  wire  GEN_2402;
  wire  GEN_2403;
  wire  GEN_2404;
  wire  GEN_2405;
  wire  GEN_2406;
  wire  GEN_2407;
  wire  GEN_2408;
  wire  GEN_2409;
  wire  GEN_2410;
  wire  GEN_2411;
  wire  GEN_2412;
  wire  GEN_2413;
  wire  GEN_2414;
  wire  GEN_2415;
  wire  GEN_2416;
  wire  GEN_2417;
  wire  GEN_2418;
  wire  GEN_2419;
  wire  GEN_2420;
  wire  GEN_2421;
  wire  GEN_2422;
  wire  GEN_2423;
  wire  GEN_2424;
  wire  GEN_2425;
  wire  GEN_2426;
  wire  GEN_2427;
  wire  GEN_2428;
  wire  GEN_2429;
  wire  GEN_2430;
  wire  GEN_2431;
  wire  GEN_2432;
  wire  GEN_2433;
  wire  GEN_2434;
  wire  GEN_2435;
  wire  GEN_2436;
  wire  GEN_2437;
  wire  GEN_2438;
  wire  GEN_2439;
  wire  GEN_2440;
  wire  GEN_2441;
  wire  GEN_2442;
  wire  GEN_2443;
  wire  GEN_2444;
  wire  GEN_2445;
  wire  GEN_2446;
  wire  GEN_2447;
  wire  GEN_2448;
  wire  GEN_2449;
  wire  GEN_2450;
  wire  GEN_2451;
  wire  GEN_2452;
  wire  GEN_2453;
  wire  GEN_2454;
  wire  GEN_2455;
  wire  GEN_2456;
  wire  GEN_2457;
  wire  GEN_2458;
  wire  GEN_2459;
  wire  GEN_2460;
  wire  GEN_2461;
  wire  GEN_2462;
  wire  GEN_2463;
  wire  GEN_2464;
  wire  GEN_2465;
  wire  GEN_2466;
  wire  T_24260;
  wire  T_24261;
  wire  T_24262;
  wire  T_24263;
  wire  T_24264;
  wire [511:0] T_24266;
  wire  T_25293;
  wire  T_25294;
  wire  T_25295;
  wire  T_25296;
  wire  T_25299;
  wire  T_25300;
  wire  T_25302;
  wire  T_25303;
  wire  T_25304;
  wire  T_25306;
  wire  T_25310;
  wire  T_25312;
  wire  T_25315;
  wire  T_25316;
  wire  T_25322;
  wire  T_25326;
  wire  T_25332;
  wire  T_25335;
  wire  T_25336;
  wire  T_25342;
  wire  T_25346;
  wire  T_25352;
  wire  T_25355;
  wire  T_25356;
  wire  T_25362;
  wire  T_25366;
  wire  T_25372;
  wire  T_25375;
  wire  T_25376;
  wire  T_25382;
  wire  T_25386;
  wire  T_25392;
  wire  T_25395;
  wire  T_25396;
  wire  T_25402;
  wire  T_25406;
  wire  T_25412;
  wire  T_25415;
  wire  T_25416;
  wire  T_25422;
  wire  T_25426;
  wire  T_25432;
  wire  T_25435;
  wire  T_25436;
  wire  T_25442;
  wire  T_25446;
  wire  T_25452;
  wire  T_25455;
  wire  T_25456;
  wire  T_25462;
  wire  T_25466;
  wire  T_25472;
  wire  T_25475;
  wire  T_25476;
  wire  T_25482;
  wire  T_25486;
  wire  T_25492;
  wire  T_25495;
  wire  T_25496;
  wire  T_25502;
  wire  T_25506;
  wire  T_25512;
  wire  T_25515;
  wire  T_25516;
  wire  T_25522;
  wire  T_25526;
  wire  T_25532;
  wire  T_25535;
  wire  T_25536;
  wire  T_25542;
  wire  T_25546;
  wire  T_25552;
  wire  T_25555;
  wire  T_25556;
  wire  T_25562;
  wire  T_25566;
  wire  T_25572;
  wire  T_25575;
  wire  T_25576;
  wire  T_25582;
  wire  T_25586;
  wire  T_25592;
  wire  T_25595;
  wire  T_25596;
  wire  T_25602;
  wire  T_25606;
  wire  T_25612;
  wire  T_25615;
  wire  T_25616;
  wire  T_25622;
  wire  T_25626;
  wire  T_25632;
  wire  T_25635;
  wire  T_25636;
  wire  T_25642;
  wire  T_25646;
  wire  T_25652;
  wire  T_25655;
  wire  T_25656;
  wire  T_25662;
  wire  T_25666;
  wire  T_25672;
  wire  T_25675;
  wire  T_25676;
  wire  T_25682;
  wire  T_25686;
  wire  T_25692;
  wire  T_25695;
  wire  T_25696;
  wire  T_25702;
  wire  T_25706;
  wire  T_25712;
  wire  T_25715;
  wire  T_25716;
  wire  T_25722;
  wire  T_25726;
  wire  T_25732;
  wire  T_25735;
  wire  T_25736;
  wire  T_25742;
  wire  T_25746;
  wire  T_25752;
  wire  T_25755;
  wire  T_25756;
  wire  T_25762;
  wire  T_25766;
  wire  T_25772;
  wire  T_25775;
  wire  T_25776;
  wire  T_25782;
  wire  T_25786;
  wire  T_25792;
  wire  T_25795;
  wire  T_25796;
  wire  T_25802;
  wire  T_25806;
  wire  T_25812;
  wire  T_25815;
  wire  T_25816;
  wire  T_25822;
  wire  T_25826;
  wire  T_25832;
  wire  T_25835;
  wire  T_25836;
  wire  T_25842;
  wire  T_25846;
  wire  T_25852;
  wire  T_25855;
  wire  T_25856;
  wire  T_25862;
  wire  T_25866;
  wire  T_25872;
  wire  T_25875;
  wire  T_25876;
  wire  T_25882;
  wire  T_25886;
  wire  T_25892;
  wire  T_25895;
  wire  T_25896;
  wire  T_25902;
  wire  T_25906;
  wire  T_25912;
  wire  T_25915;
  wire  T_25916;
  wire  T_25922;
  wire  T_25926;
  wire  T_25932;
  wire  T_25935;
  wire  T_25936;
  wire  T_25942;
  wire  T_25946;
  wire  T_25952;
  wire  T_25955;
  wire  T_25956;
  wire  T_25962;
  wire  T_25966;
  wire  T_25972;
  wire  T_25975;
  wire  T_25976;
  wire  T_25982;
  wire  T_25986;
  wire  T_25992;
  wire  T_25995;
  wire  T_25996;
  wire  T_26002;
  wire  T_26006;
  wire  T_26012;
  wire  T_26015;
  wire  T_26016;
  wire  T_26022;
  wire  T_26026;
  wire  T_26032;
  wire  T_26035;
  wire  T_26036;
  wire  T_26042;
  wire  T_26046;
  wire  T_26052;
  wire  T_26055;
  wire  T_26056;
  wire  T_26062;
  wire  T_26066;
  wire  T_26072;
  wire  T_26075;
  wire  T_26076;
  wire  T_26082;
  wire  T_26086;
  wire  T_26092;
  wire  T_26095;
  wire  T_26096;
  wire  T_26102;
  wire  T_26106;
  wire  T_26112;
  wire  T_26115;
  wire  T_26116;
  wire  T_26122;
  wire  T_26126;
  wire  T_26132;
  wire  T_26135;
  wire  T_26136;
  wire  T_26142;
  wire  T_26146;
  wire  T_26152;
  wire  T_26155;
  wire  T_26156;
  wire  T_26162;
  wire  T_26166;
  wire  T_26172;
  wire  T_26175;
  wire  T_26176;
  wire  T_26182;
  wire  T_26186;
  wire  T_26192;
  wire  T_26195;
  wire  T_26196;
  wire  T_26202;
  wire  T_26206;
  wire  T_26212;
  wire  T_26215;
  wire  T_26216;
  wire  T_26222;
  wire  T_26226;
  wire  T_26232;
  wire  T_26235;
  wire  T_26236;
  wire  T_26242;
  wire  T_26246;
  wire  T_26252;
  wire  T_26255;
  wire  T_26256;
  wire  T_26262;
  wire  T_26266;
  wire  T_26272;
  wire  T_26275;
  wire  T_26276;
  wire  T_26282;
  wire  T_26286;
  wire  T_26292;
  wire  T_26295;
  wire  T_26296;
  wire  T_26302;
  wire  T_26306;
  wire  T_26312;
  wire  T_26315;
  wire  T_26316;
  wire  T_26322;
  wire  T_26326;
  wire  T_26332;
  wire  T_26575;
  wire  T_26576;
  wire  T_26582;
  wire  T_26586;
  wire  T_26592;
  wire  T_26595;
  wire  T_26596;
  wire  T_26602;
  wire  T_26606;
  wire  T_26612;
  wire  T_27855;
  wire  T_27856;
  wire  T_27862;
  wire  T_27866;
  wire  T_27872;
  wire  T_27875;
  wire  T_27876;
  wire  T_27882;
  wire  T_27886;
  wire  T_27892;
  wire  T_30415;
  wire  T_30416;
  wire  T_30422;
  wire  T_30426;
  wire  T_30432;
  wire  T_30435;
  wire  T_30436;
  wire  T_30442;
  wire  T_30446;
  wire  T_30452;
  wire  T_35533;
  wire  T_35534;
  wire  T_35535;
  wire  T_35536;
  wire  T_35537;
  wire  T_35538;
  wire  T_35539;
  wire  T_35540;
  wire  T_35541;
  wire  T_35542;
  wire  T_35543;
  wire  T_35544;
  wire  T_35545;
  wire  T_35546;
  wire  T_35547;
  wire  T_35548;
  wire  T_35549;
  wire  T_35550;
  wire  T_35551;
  wire  T_35552;
  wire  T_35553;
  wire  T_35554;
  wire  T_35555;
  wire  T_35556;
  wire  T_35557;
  wire  T_35558;
  wire  T_35559;
  wire  T_35560;
  wire  T_35561;
  wire  T_35562;
  wire  T_35563;
  wire  T_35565;
  wire  T_35566;
  wire  T_35567;
  wire  T_35568;
  wire  T_35569;
  wire  T_35570;
  wire  T_35571;
  wire  T_35572;
  wire  T_35573;
  wire  T_35574;
  wire  T_35575;
  wire  T_35576;
  wire  T_35577;
  wire  T_35578;
  wire  T_35579;
  wire  T_35580;
  wire  T_35581;
  wire  T_35582;
  wire  T_35583;
  wire  T_35584;
  wire  T_35585;
  wire  T_35586;
  wire  T_35587;
  wire  T_35588;
  wire  T_35589;
  wire  T_35590;
  wire  T_35591;
  wire  T_35592;
  wire  T_35593;
  wire  T_35594;
  wire  T_35595;
  wire  T_35597;
  wire  T_35598;
  wire  T_35599;
  wire  T_35600;
  wire  T_35601;
  wire  T_35602;
  wire  T_35603;
  wire  T_35604;
  wire  T_35605;
  wire  T_35606;
  wire  T_35607;
  wire  T_35608;
  wire  T_35609;
  wire  T_35610;
  wire  T_35611;
  wire  T_35612;
  wire  T_35613;
  wire  T_35614;
  wire  T_35615;
  wire  T_35616;
  wire  T_35617;
  wire  T_35618;
  wire  T_35619;
  wire  T_35620;
  wire  T_35621;
  wire  T_35622;
  wire  T_35623;
  wire  T_35624;
  wire  T_35625;
  wire  T_35626;
  wire  T_35627;
  wire  T_35629;
  wire  T_35630;
  wire  T_35631;
  wire  T_35632;
  wire  T_35633;
  wire  T_35634;
  wire  T_35635;
  wire  T_35636;
  wire  T_35637;
  wire  T_35638;
  wire  T_35639;
  wire  T_35640;
  wire  T_35641;
  wire  T_35642;
  wire  T_35643;
  wire  T_35644;
  wire  T_35645;
  wire  T_35646;
  wire  T_35647;
  wire  T_35648;
  wire  T_35649;
  wire  T_35650;
  wire  T_35651;
  wire  T_35652;
  wire  T_35653;
  wire  T_35654;
  wire  T_35655;
  wire  T_35656;
  wire  T_35657;
  wire  T_35658;
  wire  T_35659;
  wire  T_35691;
  wire  T_35723;
  wire  T_35755;
  wire  T_35787;
  wire  T_35818;
  wire  T_35819;
  wire  T_35850;
  wire  T_35851;
  wire  T_35882;
  wire  T_35883;
  wire  T_35914;
  wire  T_35915;
  wire  T_35945;
  wire  T_35946;
  wire  T_35947;
  wire  T_35977;
  wire  T_35978;
  wire  T_35979;
  wire  T_36009;
  wire  T_36010;
  wire  T_36011;
  wire  T_36041;
  wire  T_36042;
  wire  T_36043;
  wire  T_36072;
  wire  T_36073;
  wire  T_36074;
  wire  T_36075;
  wire  T_36104;
  wire  T_36105;
  wire  T_36106;
  wire  T_36107;
  wire  T_36136;
  wire  T_36137;
  wire  T_36138;
  wire  T_36139;
  wire  T_36168;
  wire  T_36169;
  wire  T_36170;
  wire  T_36171;
  wire  T_36199;
  wire  T_36200;
  wire  T_36201;
  wire  T_36202;
  wire  T_36203;
  wire  T_36231;
  wire  T_36232;
  wire  T_36233;
  wire  T_36234;
  wire  T_36235;
  wire  T_36263;
  wire  T_36264;
  wire  T_36265;
  wire  T_36266;
  wire  T_36267;
  wire  T_36295;
  wire  T_36296;
  wire  T_36297;
  wire  T_36298;
  wire  T_36299;
  wire  T_36326;
  wire  T_36327;
  wire  T_36328;
  wire  T_36329;
  wire  T_36330;
  wire  T_36331;
  wire  T_36358;
  wire  T_36359;
  wire  T_36360;
  wire  T_36361;
  wire  T_36362;
  wire  T_36363;
  wire  T_36390;
  wire  T_36391;
  wire  T_36392;
  wire  T_36393;
  wire  T_36394;
  wire  T_36395;
  wire  T_36422;
  wire  T_36423;
  wire  T_36424;
  wire  T_36425;
  wire  T_36426;
  wire  T_36427;
  wire  T_36453;
  wire  T_36454;
  wire  T_36455;
  wire  T_36456;
  wire  T_36457;
  wire  T_36458;
  wire  T_36459;
  wire  T_36485;
  wire  T_36486;
  wire  T_36487;
  wire  T_36488;
  wire  T_36489;
  wire  T_36490;
  wire  T_36491;
  wire  T_36517;
  wire  T_36518;
  wire  T_36519;
  wire  T_36520;
  wire  T_36521;
  wire  T_36522;
  wire  T_36523;
  wire  T_36549;
  wire  T_36550;
  wire  T_36551;
  wire  T_36552;
  wire  T_36553;
  wire  T_36554;
  wire  T_36555;
  wire  T_36580;
  wire  T_36581;
  wire  T_36582;
  wire  T_36583;
  wire  T_36584;
  wire  T_36585;
  wire  T_36586;
  wire  T_36587;
  wire  T_36612;
  wire  T_36613;
  wire  T_36614;
  wire  T_36615;
  wire  T_36616;
  wire  T_36617;
  wire  T_36618;
  wire  T_36619;
  wire  T_36644;
  wire  T_36645;
  wire  T_36646;
  wire  T_36647;
  wire  T_36648;
  wire  T_36649;
  wire  T_36650;
  wire  T_36651;
  wire  T_36676;
  wire  T_36677;
  wire  T_36678;
  wire  T_36679;
  wire  T_36680;
  wire  T_36681;
  wire  T_36682;
  wire  T_36683;
  wire  T_36707;
  wire  T_36708;
  wire  T_36709;
  wire  T_36710;
  wire  T_36711;
  wire  T_36712;
  wire  T_36713;
  wire  T_36714;
  wire  T_36715;
  wire  T_36739;
  wire  T_36740;
  wire  T_36741;
  wire  T_36742;
  wire  T_36743;
  wire  T_36744;
  wire  T_36745;
  wire  T_36746;
  wire  T_36747;
  wire  T_36771;
  wire  T_36772;
  wire  T_36773;
  wire  T_36774;
  wire  T_36775;
  wire  T_36776;
  wire  T_36777;
  wire  T_36778;
  wire  T_36779;
  wire  T_36803;
  wire  T_36804;
  wire  T_36805;
  wire  T_36806;
  wire  T_36807;
  wire  T_36808;
  wire  T_36809;
  wire  T_36810;
  wire  T_36811;
  wire  T_36834;
  wire  T_36835;
  wire  T_36836;
  wire  T_36837;
  wire  T_36838;
  wire  T_36839;
  wire  T_36840;
  wire  T_36841;
  wire  T_36842;
  wire  T_36843;
  wire  T_36866;
  wire  T_36867;
  wire  T_36868;
  wire  T_36869;
  wire  T_36870;
  wire  T_36871;
  wire  T_36872;
  wire  T_36873;
  wire  T_36874;
  wire  T_36875;
  wire  T_36898;
  wire  T_36899;
  wire  T_36900;
  wire  T_36901;
  wire  T_36902;
  wire  T_36903;
  wire  T_36904;
  wire  T_36905;
  wire  T_36906;
  wire  T_36907;
  wire  T_36930;
  wire  T_36931;
  wire  T_36932;
  wire  T_36933;
  wire  T_36934;
  wire  T_36935;
  wire  T_36936;
  wire  T_36937;
  wire  T_36938;
  wire  T_36939;
  wire  T_36961;
  wire  T_36962;
  wire  T_36963;
  wire  T_36964;
  wire  T_36965;
  wire  T_36966;
  wire  T_36967;
  wire  T_36968;
  wire  T_36969;
  wire  T_36970;
  wire  T_36971;
  wire  T_36993;
  wire  T_36994;
  wire  T_36995;
  wire  T_36996;
  wire  T_36997;
  wire  T_36998;
  wire  T_36999;
  wire  T_37000;
  wire  T_37001;
  wire  T_37002;
  wire  T_37003;
  wire  T_37025;
  wire  T_37026;
  wire  T_37027;
  wire  T_37028;
  wire  T_37029;
  wire  T_37030;
  wire  T_37031;
  wire  T_37032;
  wire  T_37033;
  wire  T_37034;
  wire  T_37035;
  wire  T_37057;
  wire  T_37058;
  wire  T_37059;
  wire  T_37060;
  wire  T_37061;
  wire  T_37062;
  wire  T_37063;
  wire  T_37064;
  wire  T_37065;
  wire  T_37066;
  wire  T_37067;
  wire  T_37088;
  wire  T_37089;
  wire  T_37090;
  wire  T_37091;
  wire  T_37092;
  wire  T_37093;
  wire  T_37094;
  wire  T_37095;
  wire  T_37096;
  wire  T_37097;
  wire  T_37098;
  wire  T_37099;
  wire  T_37120;
  wire  T_37121;
  wire  T_37122;
  wire  T_37123;
  wire  T_37124;
  wire  T_37125;
  wire  T_37126;
  wire  T_37127;
  wire  T_37128;
  wire  T_37129;
  wire  T_37130;
  wire  T_37131;
  wire  T_37152;
  wire  T_37153;
  wire  T_37154;
  wire  T_37155;
  wire  T_37156;
  wire  T_37157;
  wire  T_37158;
  wire  T_37159;
  wire  T_37160;
  wire  T_37161;
  wire  T_37162;
  wire  T_37163;
  wire  T_37184;
  wire  T_37185;
  wire  T_37186;
  wire  T_37187;
  wire  T_37188;
  wire  T_37189;
  wire  T_37190;
  wire  T_37191;
  wire  T_37192;
  wire  T_37193;
  wire  T_37194;
  wire  T_37195;
  wire  T_37215;
  wire  T_37216;
  wire  T_37217;
  wire  T_37218;
  wire  T_37219;
  wire  T_37220;
  wire  T_37221;
  wire  T_37222;
  wire  T_37223;
  wire  T_37224;
  wire  T_37225;
  wire  T_37226;
  wire  T_37227;
  wire  T_37247;
  wire  T_37248;
  wire  T_37249;
  wire  T_37250;
  wire  T_37251;
  wire  T_37252;
  wire  T_37253;
  wire  T_37254;
  wire  T_37255;
  wire  T_37256;
  wire  T_37257;
  wire  T_37258;
  wire  T_37259;
  wire  T_37279;
  wire  T_37280;
  wire  T_37281;
  wire  T_37282;
  wire  T_37283;
  wire  T_37284;
  wire  T_37285;
  wire  T_37286;
  wire  T_37287;
  wire  T_37288;
  wire  T_37289;
  wire  T_37290;
  wire  T_37291;
  wire  T_37311;
  wire  T_37312;
  wire  T_37313;
  wire  T_37314;
  wire  T_37315;
  wire  T_37316;
  wire  T_37317;
  wire  T_37318;
  wire  T_37319;
  wire  T_37320;
  wire  T_37321;
  wire  T_37322;
  wire  T_37323;
  wire  T_37342;
  wire  T_37343;
  wire  T_37344;
  wire  T_37345;
  wire  T_37346;
  wire  T_37347;
  wire  T_37348;
  wire  T_37349;
  wire  T_37350;
  wire  T_37351;
  wire  T_37352;
  wire  T_37353;
  wire  T_37354;
  wire  T_37355;
  wire  T_37374;
  wire  T_37375;
  wire  T_37376;
  wire  T_37377;
  wire  T_37378;
  wire  T_37379;
  wire  T_37380;
  wire  T_37381;
  wire  T_37382;
  wire  T_37383;
  wire  T_37384;
  wire  T_37385;
  wire  T_37386;
  wire  T_37387;
  wire  T_37406;
  wire  T_37407;
  wire  T_37408;
  wire  T_37409;
  wire  T_37410;
  wire  T_37411;
  wire  T_37412;
  wire  T_37413;
  wire  T_37414;
  wire  T_37415;
  wire  T_37416;
  wire  T_37417;
  wire  T_37418;
  wire  T_37419;
  wire  T_37438;
  wire  T_37439;
  wire  T_37440;
  wire  T_37441;
  wire  T_37442;
  wire  T_37443;
  wire  T_37444;
  wire  T_37445;
  wire  T_37446;
  wire  T_37447;
  wire  T_37448;
  wire  T_37449;
  wire  T_37450;
  wire  T_37451;
  wire  T_37469;
  wire  T_37470;
  wire  T_37471;
  wire  T_37472;
  wire  T_37473;
  wire  T_37474;
  wire  T_37475;
  wire  T_37476;
  wire  T_37477;
  wire  T_37478;
  wire  T_37479;
  wire  T_37480;
  wire  T_37481;
  wire  T_37482;
  wire  T_37483;
  wire  T_37501;
  wire  T_37502;
  wire  T_37503;
  wire  T_37504;
  wire  T_37505;
  wire  T_37506;
  wire  T_37507;
  wire  T_37508;
  wire  T_37509;
  wire  T_37510;
  wire  T_37511;
  wire  T_37512;
  wire  T_37513;
  wire  T_37514;
  wire  T_37515;
  wire  T_37533;
  wire  T_37534;
  wire  T_37535;
  wire  T_37536;
  wire  T_37537;
  wire  T_37538;
  wire  T_37539;
  wire  T_37540;
  wire  T_37541;
  wire  T_37542;
  wire  T_37543;
  wire  T_37544;
  wire  T_37545;
  wire  T_37546;
  wire  T_37547;
  wire  T_37565;
  wire  T_37566;
  wire  T_37567;
  wire  T_37568;
  wire  T_37569;
  wire  T_37570;
  wire  T_37571;
  wire  T_37572;
  wire  T_37573;
  wire  T_37574;
  wire  T_37575;
  wire  T_37576;
  wire  T_37577;
  wire  T_37578;
  wire  T_37579;
  wire  T_37596;
  wire  T_37597;
  wire  T_37598;
  wire  T_37599;
  wire  T_37600;
  wire  T_37601;
  wire  T_37602;
  wire  T_37603;
  wire  T_37604;
  wire  T_37605;
  wire  T_37606;
  wire  T_37607;
  wire  T_37608;
  wire  T_37609;
  wire  T_37610;
  wire  T_37611;
  wire  T_37628;
  wire  T_37629;
  wire  T_37630;
  wire  T_37631;
  wire  T_37632;
  wire  T_37633;
  wire  T_37634;
  wire  T_37635;
  wire  T_37636;
  wire  T_37637;
  wire  T_37638;
  wire  T_37639;
  wire  T_37640;
  wire  T_37641;
  wire  T_37642;
  wire  T_37643;
  wire  T_37660;
  wire  T_37661;
  wire  T_37662;
  wire  T_37663;
  wire  T_37664;
  wire  T_37665;
  wire  T_37666;
  wire  T_37667;
  wire  T_37668;
  wire  T_37669;
  wire  T_37670;
  wire  T_37671;
  wire  T_37672;
  wire  T_37673;
  wire  T_37674;
  wire  T_37675;
  wire  T_37692;
  wire  T_37693;
  wire  T_37694;
  wire  T_37695;
  wire  T_37696;
  wire  T_37697;
  wire  T_37698;
  wire  T_37699;
  wire  T_37700;
  wire  T_37701;
  wire  T_37702;
  wire  T_37703;
  wire  T_37704;
  wire  T_37705;
  wire  T_37706;
  wire  T_37707;
  wire  T_37723;
  wire  T_37724;
  wire  T_37725;
  wire  T_37726;
  wire  T_37727;
  wire  T_37728;
  wire  T_37729;
  wire  T_37730;
  wire  T_37731;
  wire  T_37732;
  wire  T_37733;
  wire  T_37734;
  wire  T_37735;
  wire  T_37736;
  wire  T_37737;
  wire  T_37738;
  wire  T_37739;
  wire  T_37755;
  wire  T_37756;
  wire  T_37757;
  wire  T_37758;
  wire  T_37759;
  wire  T_37760;
  wire  T_37761;
  wire  T_37762;
  wire  T_37763;
  wire  T_37764;
  wire  T_37765;
  wire  T_37766;
  wire  T_37767;
  wire  T_37768;
  wire  T_37769;
  wire  T_37770;
  wire  T_37771;
  wire  T_37787;
  wire  T_37788;
  wire  T_37789;
  wire  T_37790;
  wire  T_37791;
  wire  T_37792;
  wire  T_37793;
  wire  T_37794;
  wire  T_37795;
  wire  T_37796;
  wire  T_37797;
  wire  T_37798;
  wire  T_37799;
  wire  T_37800;
  wire  T_37801;
  wire  T_37802;
  wire  T_37803;
  wire  T_37819;
  wire  T_37820;
  wire  T_37821;
  wire  T_37822;
  wire  T_37823;
  wire  T_37824;
  wire  T_37825;
  wire  T_37826;
  wire  T_37827;
  wire  T_37828;
  wire  T_37829;
  wire  T_37830;
  wire  T_37831;
  wire  T_37832;
  wire  T_37833;
  wire  T_37834;
  wire  T_37835;
  wire  T_37850;
  wire  T_37851;
  wire  T_37852;
  wire  T_37853;
  wire  T_37854;
  wire  T_37855;
  wire  T_37856;
  wire  T_37857;
  wire  T_37858;
  wire  T_37859;
  wire  T_37860;
  wire  T_37861;
  wire  T_37862;
  wire  T_37863;
  wire  T_37864;
  wire  T_37865;
  wire  T_37866;
  wire  T_37867;
  wire  T_37882;
  wire  T_37883;
  wire  T_37884;
  wire  T_37885;
  wire  T_37886;
  wire  T_37887;
  wire  T_37888;
  wire  T_37889;
  wire  T_37890;
  wire  T_37891;
  wire  T_37892;
  wire  T_37893;
  wire  T_37894;
  wire  T_37895;
  wire  T_37896;
  wire  T_37897;
  wire  T_37898;
  wire  T_37899;
  wire  T_37914;
  wire  T_37915;
  wire  T_37916;
  wire  T_37917;
  wire  T_37918;
  wire  T_37919;
  wire  T_37920;
  wire  T_37921;
  wire  T_37922;
  wire  T_37923;
  wire  T_37924;
  wire  T_37925;
  wire  T_37926;
  wire  T_37927;
  wire  T_37928;
  wire  T_37929;
  wire  T_37930;
  wire  T_37931;
  wire  T_37946;
  wire  T_37947;
  wire  T_37948;
  wire  T_37949;
  wire  T_37950;
  wire  T_37951;
  wire  T_37952;
  wire  T_37953;
  wire  T_37954;
  wire  T_37955;
  wire  T_37956;
  wire  T_37957;
  wire  T_37958;
  wire  T_37959;
  wire  T_37960;
  wire  T_37961;
  wire  T_37962;
  wire  T_37963;
  wire  T_37977;
  wire  T_37978;
  wire  T_37979;
  wire  T_37980;
  wire  T_37981;
  wire  T_37982;
  wire  T_37983;
  wire  T_37984;
  wire  T_37985;
  wire  T_37986;
  wire  T_37987;
  wire  T_37988;
  wire  T_37989;
  wire  T_37990;
  wire  T_37991;
  wire  T_37992;
  wire  T_37993;
  wire  T_37994;
  wire  T_37995;
  wire  T_38009;
  wire  T_38010;
  wire  T_38011;
  wire  T_38012;
  wire  T_38013;
  wire  T_38014;
  wire  T_38015;
  wire  T_38016;
  wire  T_38017;
  wire  T_38018;
  wire  T_38019;
  wire  T_38020;
  wire  T_38021;
  wire  T_38022;
  wire  T_38023;
  wire  T_38024;
  wire  T_38025;
  wire  T_38026;
  wire  T_38027;
  wire  T_38041;
  wire  T_38042;
  wire  T_38043;
  wire  T_38044;
  wire  T_38045;
  wire  T_38046;
  wire  T_38047;
  wire  T_38048;
  wire  T_38049;
  wire  T_38050;
  wire  T_38051;
  wire  T_38052;
  wire  T_38053;
  wire  T_38054;
  wire  T_38055;
  wire  T_38056;
  wire  T_38057;
  wire  T_38058;
  wire  T_38059;
  wire  T_38073;
  wire  T_38074;
  wire  T_38075;
  wire  T_38076;
  wire  T_38077;
  wire  T_38078;
  wire  T_38079;
  wire  T_38080;
  wire  T_38081;
  wire  T_38082;
  wire  T_38083;
  wire  T_38084;
  wire  T_38085;
  wire  T_38086;
  wire  T_38087;
  wire  T_38088;
  wire  T_38089;
  wire  T_38090;
  wire  T_38091;
  wire  T_38104;
  wire  T_38105;
  wire  T_38106;
  wire  T_38107;
  wire  T_38108;
  wire  T_38109;
  wire  T_38110;
  wire  T_38111;
  wire  T_38112;
  wire  T_38113;
  wire  T_38114;
  wire  T_38115;
  wire  T_38116;
  wire  T_38117;
  wire  T_38118;
  wire  T_38119;
  wire  T_38120;
  wire  T_38121;
  wire  T_38122;
  wire  T_38123;
  wire  T_38136;
  wire  T_38137;
  wire  T_38138;
  wire  T_38139;
  wire  T_38140;
  wire  T_38141;
  wire  T_38142;
  wire  T_38143;
  wire  T_38144;
  wire  T_38145;
  wire  T_38146;
  wire  T_38147;
  wire  T_38148;
  wire  T_38149;
  wire  T_38150;
  wire  T_38151;
  wire  T_38152;
  wire  T_38153;
  wire  T_38154;
  wire  T_38155;
  wire  T_38168;
  wire  T_38169;
  wire  T_38170;
  wire  T_38171;
  wire  T_38172;
  wire  T_38173;
  wire  T_38174;
  wire  T_38175;
  wire  T_38176;
  wire  T_38177;
  wire  T_38178;
  wire  T_38179;
  wire  T_38180;
  wire  T_38181;
  wire  T_38182;
  wire  T_38183;
  wire  T_38184;
  wire  T_38185;
  wire  T_38186;
  wire  T_38187;
  wire  T_38200;
  wire  T_38201;
  wire  T_38202;
  wire  T_38203;
  wire  T_38204;
  wire  T_38205;
  wire  T_38206;
  wire  T_38207;
  wire  T_38208;
  wire  T_38209;
  wire  T_38210;
  wire  T_38211;
  wire  T_38212;
  wire  T_38213;
  wire  T_38214;
  wire  T_38215;
  wire  T_38216;
  wire  T_38217;
  wire  T_38218;
  wire  T_38219;
  wire  T_38231;
  wire  T_38232;
  wire  T_38233;
  wire  T_38234;
  wire  T_38235;
  wire  T_38236;
  wire  T_38237;
  wire  T_38238;
  wire  T_38239;
  wire  T_38240;
  wire  T_38241;
  wire  T_38242;
  wire  T_38243;
  wire  T_38244;
  wire  T_38245;
  wire  T_38246;
  wire  T_38247;
  wire  T_38248;
  wire  T_38249;
  wire  T_38250;
  wire  T_38251;
  wire  T_38263;
  wire  T_38264;
  wire  T_38265;
  wire  T_38266;
  wire  T_38267;
  wire  T_38268;
  wire  T_38269;
  wire  T_38270;
  wire  T_38271;
  wire  T_38272;
  wire  T_38273;
  wire  T_38274;
  wire  T_38275;
  wire  T_38276;
  wire  T_38277;
  wire  T_38278;
  wire  T_38279;
  wire  T_38280;
  wire  T_38281;
  wire  T_38282;
  wire  T_38283;
  wire  T_38295;
  wire  T_38296;
  wire  T_38297;
  wire  T_38298;
  wire  T_38299;
  wire  T_38300;
  wire  T_38301;
  wire  T_38302;
  wire  T_38303;
  wire  T_38304;
  wire  T_38305;
  wire  T_38306;
  wire  T_38307;
  wire  T_38308;
  wire  T_38309;
  wire  T_38310;
  wire  T_38311;
  wire  T_38312;
  wire  T_38313;
  wire  T_38314;
  wire  T_38315;
  wire  T_38327;
  wire  T_38328;
  wire  T_38329;
  wire  T_38330;
  wire  T_38331;
  wire  T_38332;
  wire  T_38333;
  wire  T_38334;
  wire  T_38335;
  wire  T_38336;
  wire  T_38337;
  wire  T_38338;
  wire  T_38339;
  wire  T_38340;
  wire  T_38341;
  wire  T_38342;
  wire  T_38343;
  wire  T_38344;
  wire  T_38345;
  wire  T_38346;
  wire  T_38347;
  wire  T_38358;
  wire  T_38359;
  wire  T_38360;
  wire  T_38361;
  wire  T_38362;
  wire  T_38363;
  wire  T_38364;
  wire  T_38365;
  wire  T_38366;
  wire  T_38367;
  wire  T_38368;
  wire  T_38369;
  wire  T_38370;
  wire  T_38371;
  wire  T_38372;
  wire  T_38373;
  wire  T_38374;
  wire  T_38375;
  wire  T_38376;
  wire  T_38377;
  wire  T_38378;
  wire  T_38379;
  wire  T_38390;
  wire  T_38391;
  wire  T_38392;
  wire  T_38393;
  wire  T_38394;
  wire  T_38395;
  wire  T_38396;
  wire  T_38397;
  wire  T_38398;
  wire  T_38399;
  wire  T_38400;
  wire  T_38401;
  wire  T_38402;
  wire  T_38403;
  wire  T_38404;
  wire  T_38405;
  wire  T_38406;
  wire  T_38407;
  wire  T_38408;
  wire  T_38409;
  wire  T_38410;
  wire  T_38411;
  wire  T_38422;
  wire  T_38423;
  wire  T_38424;
  wire  T_38425;
  wire  T_38426;
  wire  T_38427;
  wire  T_38428;
  wire  T_38429;
  wire  T_38430;
  wire  T_38431;
  wire  T_38432;
  wire  T_38433;
  wire  T_38434;
  wire  T_38435;
  wire  T_38436;
  wire  T_38437;
  wire  T_38438;
  wire  T_38439;
  wire  T_38440;
  wire  T_38441;
  wire  T_38442;
  wire  T_38443;
  wire  T_38454;
  wire  T_38455;
  wire  T_38456;
  wire  T_38457;
  wire  T_38458;
  wire  T_38459;
  wire  T_38460;
  wire  T_38461;
  wire  T_38462;
  wire  T_38463;
  wire  T_38464;
  wire  T_38465;
  wire  T_38466;
  wire  T_38467;
  wire  T_38468;
  wire  T_38469;
  wire  T_38470;
  wire  T_38471;
  wire  T_38472;
  wire  T_38473;
  wire  T_38474;
  wire  T_38475;
  wire  T_38485;
  wire  T_38486;
  wire  T_38487;
  wire  T_38488;
  wire  T_38489;
  wire  T_38490;
  wire  T_38491;
  wire  T_38492;
  wire  T_38493;
  wire  T_38494;
  wire  T_38495;
  wire  T_38496;
  wire  T_38497;
  wire  T_38498;
  wire  T_38499;
  wire  T_38500;
  wire  T_38501;
  wire  T_38502;
  wire  T_38503;
  wire  T_38504;
  wire  T_38505;
  wire  T_38506;
  wire  T_38507;
  wire  T_38517;
  wire  T_38518;
  wire  T_38519;
  wire  T_38520;
  wire  T_38521;
  wire  T_38522;
  wire  T_38523;
  wire  T_38524;
  wire  T_38525;
  wire  T_38526;
  wire  T_38527;
  wire  T_38528;
  wire  T_38529;
  wire  T_38530;
  wire  T_38531;
  wire  T_38532;
  wire  T_38533;
  wire  T_38534;
  wire  T_38535;
  wire  T_38536;
  wire  T_38537;
  wire  T_38538;
  wire  T_38539;
  wire  T_38549;
  wire  T_38550;
  wire  T_38551;
  wire  T_38552;
  wire  T_38553;
  wire  T_38554;
  wire  T_38555;
  wire  T_38556;
  wire  T_38557;
  wire  T_38558;
  wire  T_38559;
  wire  T_38560;
  wire  T_38561;
  wire  T_38562;
  wire  T_38563;
  wire  T_38564;
  wire  T_38565;
  wire  T_38566;
  wire  T_38567;
  wire  T_38568;
  wire  T_38569;
  wire  T_38570;
  wire  T_38571;
  wire  T_38581;
  wire  T_38582;
  wire  T_38583;
  wire  T_38584;
  wire  T_38585;
  wire  T_38586;
  wire  T_38587;
  wire  T_38588;
  wire  T_38589;
  wire  T_38590;
  wire  T_38591;
  wire  T_38592;
  wire  T_38593;
  wire  T_38594;
  wire  T_38595;
  wire  T_38596;
  wire  T_38597;
  wire  T_38598;
  wire  T_38599;
  wire  T_38600;
  wire  T_38601;
  wire  T_38602;
  wire  T_38603;
  wire  T_38612;
  wire  T_38613;
  wire  T_38614;
  wire  T_38615;
  wire  T_38616;
  wire  T_38617;
  wire  T_38618;
  wire  T_38619;
  wire  T_38620;
  wire  T_38621;
  wire  T_38622;
  wire  T_38623;
  wire  T_38624;
  wire  T_38625;
  wire  T_38626;
  wire  T_38627;
  wire  T_38628;
  wire  T_38629;
  wire  T_38630;
  wire  T_38631;
  wire  T_38632;
  wire  T_38633;
  wire  T_38634;
  wire  T_38635;
  wire  T_38644;
  wire  T_38645;
  wire  T_38646;
  wire  T_38647;
  wire  T_38648;
  wire  T_38649;
  wire  T_38650;
  wire  T_38651;
  wire  T_38652;
  wire  T_38653;
  wire  T_38654;
  wire  T_38655;
  wire  T_38656;
  wire  T_38657;
  wire  T_38658;
  wire  T_38659;
  wire  T_38660;
  wire  T_38661;
  wire  T_38662;
  wire  T_38663;
  wire  T_38664;
  wire  T_38665;
  wire  T_38666;
  wire  T_38667;
  wire  T_38676;
  wire  T_38677;
  wire  T_38678;
  wire  T_38679;
  wire  T_38680;
  wire  T_38681;
  wire  T_38682;
  wire  T_38683;
  wire  T_38684;
  wire  T_38685;
  wire  T_38686;
  wire  T_38687;
  wire  T_38688;
  wire  T_38689;
  wire  T_38690;
  wire  T_38691;
  wire  T_38692;
  wire  T_38693;
  wire  T_38694;
  wire  T_38695;
  wire  T_38696;
  wire  T_38697;
  wire  T_38698;
  wire  T_38699;
  wire  T_38708;
  wire  T_38709;
  wire  T_38710;
  wire  T_38711;
  wire  T_38712;
  wire  T_38713;
  wire  T_38714;
  wire  T_38715;
  wire  T_38716;
  wire  T_38717;
  wire  T_38718;
  wire  T_38719;
  wire  T_38720;
  wire  T_38721;
  wire  T_38722;
  wire  T_38723;
  wire  T_38724;
  wire  T_38725;
  wire  T_38726;
  wire  T_38727;
  wire  T_38728;
  wire  T_38729;
  wire  T_38730;
  wire  T_38731;
  wire  T_38739;
  wire  T_38740;
  wire  T_38741;
  wire  T_38742;
  wire  T_38743;
  wire  T_38744;
  wire  T_38745;
  wire  T_38746;
  wire  T_38747;
  wire  T_38748;
  wire  T_38749;
  wire  T_38750;
  wire  T_38751;
  wire  T_38752;
  wire  T_38753;
  wire  T_38754;
  wire  T_38755;
  wire  T_38756;
  wire  T_38757;
  wire  T_38758;
  wire  T_38759;
  wire  T_38760;
  wire  T_38761;
  wire  T_38762;
  wire  T_38763;
  wire  T_38771;
  wire  T_38772;
  wire  T_38773;
  wire  T_38774;
  wire  T_38775;
  wire  T_38776;
  wire  T_38777;
  wire  T_38778;
  wire  T_38779;
  wire  T_38780;
  wire  T_38781;
  wire  T_38782;
  wire  T_38783;
  wire  T_38784;
  wire  T_38785;
  wire  T_38786;
  wire  T_38787;
  wire  T_38788;
  wire  T_38789;
  wire  T_38790;
  wire  T_38791;
  wire  T_38792;
  wire  T_38793;
  wire  T_38794;
  wire  T_38795;
  wire  T_38803;
  wire  T_38804;
  wire  T_38805;
  wire  T_38806;
  wire  T_38807;
  wire  T_38808;
  wire  T_38809;
  wire  T_38810;
  wire  T_38811;
  wire  T_38812;
  wire  T_38813;
  wire  T_38814;
  wire  T_38815;
  wire  T_38816;
  wire  T_38817;
  wire  T_38818;
  wire  T_38819;
  wire  T_38820;
  wire  T_38821;
  wire  T_38822;
  wire  T_38823;
  wire  T_38824;
  wire  T_38825;
  wire  T_38826;
  wire  T_38827;
  wire  T_38835;
  wire  T_38836;
  wire  T_38837;
  wire  T_38838;
  wire  T_38839;
  wire  T_38840;
  wire  T_38841;
  wire  T_38842;
  wire  T_38843;
  wire  T_38844;
  wire  T_38845;
  wire  T_38846;
  wire  T_38847;
  wire  T_38848;
  wire  T_38849;
  wire  T_38850;
  wire  T_38851;
  wire  T_38852;
  wire  T_38853;
  wire  T_38854;
  wire  T_38855;
  wire  T_38856;
  wire  T_38857;
  wire  T_38858;
  wire  T_38859;
  wire  T_38866;
  wire  T_38867;
  wire  T_38868;
  wire  T_38869;
  wire  T_38870;
  wire  T_38871;
  wire  T_38872;
  wire  T_38873;
  wire  T_38874;
  wire  T_38875;
  wire  T_38876;
  wire  T_38877;
  wire  T_38878;
  wire  T_38879;
  wire  T_38880;
  wire  T_38881;
  wire  T_38882;
  wire  T_38883;
  wire  T_38884;
  wire  T_38885;
  wire  T_38886;
  wire  T_38887;
  wire  T_38888;
  wire  T_38889;
  wire  T_38890;
  wire  T_38891;
  wire  T_38898;
  wire  T_38899;
  wire  T_38900;
  wire  T_38901;
  wire  T_38902;
  wire  T_38903;
  wire  T_38904;
  wire  T_38905;
  wire  T_38906;
  wire  T_38907;
  wire  T_38908;
  wire  T_38909;
  wire  T_38910;
  wire  T_38911;
  wire  T_38912;
  wire  T_38913;
  wire  T_38914;
  wire  T_38915;
  wire  T_38916;
  wire  T_38917;
  wire  T_38918;
  wire  T_38919;
  wire  T_38920;
  wire  T_38921;
  wire  T_38922;
  wire  T_38923;
  wire  T_38930;
  wire  T_38931;
  wire  T_38932;
  wire  T_38933;
  wire  T_38934;
  wire  T_38935;
  wire  T_38936;
  wire  T_38937;
  wire  T_38938;
  wire  T_38939;
  wire  T_38940;
  wire  T_38941;
  wire  T_38942;
  wire  T_38943;
  wire  T_38944;
  wire  T_38945;
  wire  T_38946;
  wire  T_38947;
  wire  T_38948;
  wire  T_38949;
  wire  T_38950;
  wire  T_38951;
  wire  T_38952;
  wire  T_38953;
  wire  T_38954;
  wire  T_38955;
  wire  T_38962;
  wire  T_38963;
  wire  T_38964;
  wire  T_38965;
  wire  T_38966;
  wire  T_38967;
  wire  T_38968;
  wire  T_38969;
  wire  T_38970;
  wire  T_38971;
  wire  T_38972;
  wire  T_38973;
  wire  T_38974;
  wire  T_38975;
  wire  T_38976;
  wire  T_38977;
  wire  T_38978;
  wire  T_38979;
  wire  T_38980;
  wire  T_38981;
  wire  T_38982;
  wire  T_38983;
  wire  T_38984;
  wire  T_38985;
  wire  T_38986;
  wire  T_38987;
  wire  T_38993;
  wire  T_38994;
  wire  T_38995;
  wire  T_38996;
  wire  T_38997;
  wire  T_38998;
  wire  T_38999;
  wire  T_39000;
  wire  T_39001;
  wire  T_39002;
  wire  T_39003;
  wire  T_39004;
  wire  T_39005;
  wire  T_39006;
  wire  T_39007;
  wire  T_39008;
  wire  T_39009;
  wire  T_39010;
  wire  T_39011;
  wire  T_39012;
  wire  T_39013;
  wire  T_39014;
  wire  T_39015;
  wire  T_39016;
  wire  T_39017;
  wire  T_39018;
  wire  T_39019;
  wire  T_39025;
  wire  T_39026;
  wire  T_39027;
  wire  T_39028;
  wire  T_39029;
  wire  T_39030;
  wire  T_39031;
  wire  T_39032;
  wire  T_39033;
  wire  T_39034;
  wire  T_39035;
  wire  T_39036;
  wire  T_39037;
  wire  T_39038;
  wire  T_39039;
  wire  T_39040;
  wire  T_39041;
  wire  T_39042;
  wire  T_39043;
  wire  T_39044;
  wire  T_39045;
  wire  T_39046;
  wire  T_39047;
  wire  T_39048;
  wire  T_39049;
  wire  T_39050;
  wire  T_39051;
  wire  T_39057;
  wire  T_39058;
  wire  T_39059;
  wire  T_39060;
  wire  T_39061;
  wire  T_39062;
  wire  T_39063;
  wire  T_39064;
  wire  T_39065;
  wire  T_39066;
  wire  T_39067;
  wire  T_39068;
  wire  T_39069;
  wire  T_39070;
  wire  T_39071;
  wire  T_39072;
  wire  T_39073;
  wire  T_39074;
  wire  T_39075;
  wire  T_39076;
  wire  T_39077;
  wire  T_39078;
  wire  T_39079;
  wire  T_39080;
  wire  T_39081;
  wire  T_39082;
  wire  T_39083;
  wire  T_39089;
  wire  T_39090;
  wire  T_39091;
  wire  T_39092;
  wire  T_39093;
  wire  T_39094;
  wire  T_39095;
  wire  T_39096;
  wire  T_39097;
  wire  T_39098;
  wire  T_39099;
  wire  T_39100;
  wire  T_39101;
  wire  T_39102;
  wire  T_39103;
  wire  T_39104;
  wire  T_39105;
  wire  T_39106;
  wire  T_39107;
  wire  T_39108;
  wire  T_39109;
  wire  T_39110;
  wire  T_39111;
  wire  T_39112;
  wire  T_39113;
  wire  T_39114;
  wire  T_39115;
  wire  T_39120;
  wire  T_39121;
  wire  T_39122;
  wire  T_39123;
  wire  T_39124;
  wire  T_39125;
  wire  T_39126;
  wire  T_39127;
  wire  T_39128;
  wire  T_39129;
  wire  T_39130;
  wire  T_39131;
  wire  T_39132;
  wire  T_39133;
  wire  T_39134;
  wire  T_39135;
  wire  T_39136;
  wire  T_39137;
  wire  T_39138;
  wire  T_39139;
  wire  T_39140;
  wire  T_39141;
  wire  T_39142;
  wire  T_39143;
  wire  T_39144;
  wire  T_39145;
  wire  T_39146;
  wire  T_39147;
  wire  T_39152;
  wire  T_39153;
  wire  T_39154;
  wire  T_39155;
  wire  T_39156;
  wire  T_39157;
  wire  T_39158;
  wire  T_39159;
  wire  T_39160;
  wire  T_39161;
  wire  T_39162;
  wire  T_39163;
  wire  T_39164;
  wire  T_39165;
  wire  T_39166;
  wire  T_39167;
  wire  T_39168;
  wire  T_39169;
  wire  T_39170;
  wire  T_39171;
  wire  T_39172;
  wire  T_39173;
  wire  T_39174;
  wire  T_39175;
  wire  T_39176;
  wire  T_39177;
  wire  T_39178;
  wire  T_39179;
  wire  T_39184;
  wire  T_39185;
  wire  T_39186;
  wire  T_39187;
  wire  T_39188;
  wire  T_39189;
  wire  T_39190;
  wire  T_39191;
  wire  T_39192;
  wire  T_39193;
  wire  T_39194;
  wire  T_39195;
  wire  T_39196;
  wire  T_39197;
  wire  T_39198;
  wire  T_39199;
  wire  T_39200;
  wire  T_39201;
  wire  T_39202;
  wire  T_39203;
  wire  T_39204;
  wire  T_39205;
  wire  T_39206;
  wire  T_39207;
  wire  T_39208;
  wire  T_39209;
  wire  T_39210;
  wire  T_39211;
  wire  T_39216;
  wire  T_39217;
  wire  T_39218;
  wire  T_39219;
  wire  T_39220;
  wire  T_39221;
  wire  T_39222;
  wire  T_39223;
  wire  T_39224;
  wire  T_39225;
  wire  T_39226;
  wire  T_39227;
  wire  T_39228;
  wire  T_39229;
  wire  T_39230;
  wire  T_39231;
  wire  T_39232;
  wire  T_39233;
  wire  T_39234;
  wire  T_39235;
  wire  T_39236;
  wire  T_39237;
  wire  T_39238;
  wire  T_39239;
  wire  T_39240;
  wire  T_39241;
  wire  T_39242;
  wire  T_39243;
  wire  T_39247;
  wire  T_39248;
  wire  T_39249;
  wire  T_39250;
  wire  T_39251;
  wire  T_39252;
  wire  T_39253;
  wire  T_39254;
  wire  T_39255;
  wire  T_39256;
  wire  T_39257;
  wire  T_39258;
  wire  T_39259;
  wire  T_39260;
  wire  T_39261;
  wire  T_39262;
  wire  T_39263;
  wire  T_39264;
  wire  T_39265;
  wire  T_39266;
  wire  T_39267;
  wire  T_39268;
  wire  T_39269;
  wire  T_39270;
  wire  T_39271;
  wire  T_39272;
  wire  T_39273;
  wire  T_39274;
  wire  T_39275;
  wire  T_39279;
  wire  T_39280;
  wire  T_39281;
  wire  T_39282;
  wire  T_39283;
  wire  T_39284;
  wire  T_39285;
  wire  T_39286;
  wire  T_39287;
  wire  T_39288;
  wire  T_39289;
  wire  T_39290;
  wire  T_39291;
  wire  T_39292;
  wire  T_39293;
  wire  T_39294;
  wire  T_39295;
  wire  T_39296;
  wire  T_39297;
  wire  T_39298;
  wire  T_39299;
  wire  T_39300;
  wire  T_39301;
  wire  T_39302;
  wire  T_39303;
  wire  T_39304;
  wire  T_39305;
  wire  T_39306;
  wire  T_39307;
  wire  T_39311;
  wire  T_39312;
  wire  T_39313;
  wire  T_39314;
  wire  T_39315;
  wire  T_39316;
  wire  T_39317;
  wire  T_39318;
  wire  T_39319;
  wire  T_39320;
  wire  T_39321;
  wire  T_39322;
  wire  T_39323;
  wire  T_39324;
  wire  T_39325;
  wire  T_39326;
  wire  T_39327;
  wire  T_39328;
  wire  T_39329;
  wire  T_39330;
  wire  T_39331;
  wire  T_39332;
  wire  T_39333;
  wire  T_39334;
  wire  T_39335;
  wire  T_39336;
  wire  T_39337;
  wire  T_39338;
  wire  T_39339;
  wire  T_39343;
  wire  T_39344;
  wire  T_39345;
  wire  T_39346;
  wire  T_39347;
  wire  T_39348;
  wire  T_39349;
  wire  T_39350;
  wire  T_39351;
  wire  T_39352;
  wire  T_39353;
  wire  T_39354;
  wire  T_39355;
  wire  T_39356;
  wire  T_39357;
  wire  T_39358;
  wire  T_39359;
  wire  T_39360;
  wire  T_39361;
  wire  T_39362;
  wire  T_39363;
  wire  T_39364;
  wire  T_39365;
  wire  T_39366;
  wire  T_39367;
  wire  T_39368;
  wire  T_39369;
  wire  T_39370;
  wire  T_39371;
  wire  T_39374;
  wire  T_39375;
  wire  T_39376;
  wire  T_39377;
  wire  T_39378;
  wire  T_39379;
  wire  T_39380;
  wire  T_39381;
  wire  T_39382;
  wire  T_39383;
  wire  T_39384;
  wire  T_39385;
  wire  T_39386;
  wire  T_39387;
  wire  T_39388;
  wire  T_39389;
  wire  T_39390;
  wire  T_39391;
  wire  T_39392;
  wire  T_39393;
  wire  T_39394;
  wire  T_39395;
  wire  T_39396;
  wire  T_39397;
  wire  T_39398;
  wire  T_39399;
  wire  T_39400;
  wire  T_39401;
  wire  T_39402;
  wire  T_39403;
  wire  T_39406;
  wire  T_39407;
  wire  T_39408;
  wire  T_39409;
  wire  T_39410;
  wire  T_39411;
  wire  T_39412;
  wire  T_39413;
  wire  T_39414;
  wire  T_39415;
  wire  T_39416;
  wire  T_39417;
  wire  T_39418;
  wire  T_39419;
  wire  T_39420;
  wire  T_39421;
  wire  T_39422;
  wire  T_39423;
  wire  T_39424;
  wire  T_39425;
  wire  T_39426;
  wire  T_39427;
  wire  T_39428;
  wire  T_39429;
  wire  T_39430;
  wire  T_39431;
  wire  T_39432;
  wire  T_39433;
  wire  T_39434;
  wire  T_39435;
  wire  T_39438;
  wire  T_39439;
  wire  T_39440;
  wire  T_39441;
  wire  T_39442;
  wire  T_39443;
  wire  T_39444;
  wire  T_39445;
  wire  T_39446;
  wire  T_39447;
  wire  T_39448;
  wire  T_39449;
  wire  T_39450;
  wire  T_39451;
  wire  T_39452;
  wire  T_39453;
  wire  T_39454;
  wire  T_39455;
  wire  T_39456;
  wire  T_39457;
  wire  T_39458;
  wire  T_39459;
  wire  T_39460;
  wire  T_39461;
  wire  T_39462;
  wire  T_39463;
  wire  T_39464;
  wire  T_39465;
  wire  T_39466;
  wire  T_39467;
  wire  T_39470;
  wire  T_39471;
  wire  T_39472;
  wire  T_39473;
  wire  T_39474;
  wire  T_39475;
  wire  T_39476;
  wire  T_39477;
  wire  T_39478;
  wire  T_39479;
  wire  T_39480;
  wire  T_39481;
  wire  T_39482;
  wire  T_39483;
  wire  T_39484;
  wire  T_39485;
  wire  T_39486;
  wire  T_39487;
  wire  T_39488;
  wire  T_39489;
  wire  T_39490;
  wire  T_39491;
  wire  T_39492;
  wire  T_39493;
  wire  T_39494;
  wire  T_39495;
  wire  T_39496;
  wire  T_39497;
  wire  T_39498;
  wire  T_39499;
  wire  T_39501;
  wire  T_39502;
  wire  T_39503;
  wire  T_39504;
  wire  T_39505;
  wire  T_39506;
  wire  T_39507;
  wire  T_39508;
  wire  T_39509;
  wire  T_39510;
  wire  T_39511;
  wire  T_39512;
  wire  T_39513;
  wire  T_39514;
  wire  T_39515;
  wire  T_39516;
  wire  T_39517;
  wire  T_39518;
  wire  T_39519;
  wire  T_39520;
  wire  T_39521;
  wire  T_39522;
  wire  T_39523;
  wire  T_39524;
  wire  T_39525;
  wire  T_39526;
  wire  T_39527;
  wire  T_39528;
  wire  T_39529;
  wire  T_39530;
  wire  T_39531;
  wire  T_39533;
  wire  T_39534;
  wire  T_39535;
  wire  T_39536;
  wire  T_39537;
  wire  T_39538;
  wire  T_39539;
  wire  T_39540;
  wire  T_39541;
  wire  T_39542;
  wire  T_39543;
  wire  T_39544;
  wire  T_39545;
  wire  T_39546;
  wire  T_39547;
  wire  T_39548;
  wire  T_39549;
  wire  T_39550;
  wire  T_39551;
  wire  T_39552;
  wire  T_39553;
  wire  T_39554;
  wire  T_39555;
  wire  T_39556;
  wire  T_39557;
  wire  T_39558;
  wire  T_39559;
  wire  T_39560;
  wire  T_39561;
  wire  T_39562;
  wire  T_39563;
  wire  T_39565;
  wire  T_39566;
  wire  T_39567;
  wire  T_39568;
  wire  T_39569;
  wire  T_39570;
  wire  T_39571;
  wire  T_39572;
  wire  T_39573;
  wire  T_39574;
  wire  T_39575;
  wire  T_39576;
  wire  T_39577;
  wire  T_39578;
  wire  T_39579;
  wire  T_39580;
  wire  T_39581;
  wire  T_39582;
  wire  T_39583;
  wire  T_39584;
  wire  T_39585;
  wire  T_39586;
  wire  T_39587;
  wire  T_39588;
  wire  T_39589;
  wire  T_39590;
  wire  T_39591;
  wire  T_39592;
  wire  T_39593;
  wire  T_39594;
  wire  T_39595;
  wire  T_39597;
  wire  T_39598;
  wire  T_39599;
  wire  T_39600;
  wire  T_39601;
  wire  T_39602;
  wire  T_39603;
  wire  T_39604;
  wire  T_39605;
  wire  T_39606;
  wire  T_39607;
  wire  T_39608;
  wire  T_39609;
  wire  T_39610;
  wire  T_39611;
  wire  T_39612;
  wire  T_39613;
  wire  T_39614;
  wire  T_39615;
  wire  T_39616;
  wire  T_39617;
  wire  T_39618;
  wire  T_39619;
  wire  T_39620;
  wire  T_39621;
  wire  T_39622;
  wire  T_39623;
  wire  T_39624;
  wire  T_39625;
  wire  T_39626;
  wire  T_39627;
  wire  T_39665;
  wire  T_39666;
  wire  T_39667;
  wire  T_39668;
  wire  T_39669;
  wire  T_39670;
  wire  T_39671;
  wire  T_39672;
  wire  T_39673;
  wire  T_39674;
  wire  T_39675;
  wire  T_39676;
  wire  T_39677;
  wire  T_39678;
  wire  T_39679;
  wire  T_39680;
  wire  T_39681;
  wire  T_39682;
  wire  T_39683;
  wire  T_39685;
  wire  T_39686;
  wire  T_39687;
  wire  T_39688;
  wire  T_39689;
  wire  T_39690;
  wire  T_39691;
  wire  T_39692;
  wire  T_39693;
  wire  T_39694;
  wire  T_39695;
  wire  T_39696;
  wire  T_39697;
  wire  T_39698;
  wire  T_39699;
  wire  T_39700;
  wire  T_39701;
  wire  T_39702;
  wire  T_39703;
  wire  T_39705;
  wire  T_39706;
  wire  T_39707;
  wire  T_39708;
  wire  T_39709;
  wire  T_39710;
  wire  T_39711;
  wire  T_39712;
  wire  T_39713;
  wire  T_39714;
  wire  T_39715;
  wire  T_39716;
  wire  T_39717;
  wire  T_39718;
  wire  T_39719;
  wire  T_39720;
  wire  T_39721;
  wire  T_39722;
  wire  T_39723;
  wire  T_39725;
  wire  T_39726;
  wire  T_39727;
  wire  T_39728;
  wire  T_39729;
  wire  T_39730;
  wire  T_39731;
  wire  T_39732;
  wire  T_39733;
  wire  T_39734;
  wire  T_39735;
  wire  T_39736;
  wire  T_39737;
  wire  T_39738;
  wire  T_39739;
  wire  T_39740;
  wire  T_39741;
  wire  T_39742;
  wire  T_39743;
  wire  T_39763;
  wire  T_39783;
  wire  T_39803;
  wire  T_39823;
  wire  T_39842;
  wire  T_39843;
  wire  T_39862;
  wire  T_39863;
  wire  T_39882;
  wire  T_39883;
  wire  T_39902;
  wire  T_39903;
  wire  T_39921;
  wire  T_39922;
  wire  T_39923;
  wire  T_39941;
  wire  T_39942;
  wire  T_39943;
  wire  T_39961;
  wire  T_39962;
  wire  T_39963;
  wire  T_39981;
  wire  T_39982;
  wire  T_39983;
  wire  T_40000;
  wire  T_40001;
  wire  T_40002;
  wire  T_40003;
  wire  T_40020;
  wire  T_40021;
  wire  T_40022;
  wire  T_40023;
  wire  T_40040;
  wire  T_40041;
  wire  T_40042;
  wire  T_40043;
  wire  T_40060;
  wire  T_40061;
  wire  T_40062;
  wire  T_40063;
  wire  T_40079;
  wire  T_40080;
  wire  T_40081;
  wire  T_40082;
  wire  T_40083;
  wire  T_40099;
  wire  T_40100;
  wire  T_40101;
  wire  T_40102;
  wire  T_40103;
  wire  T_40119;
  wire  T_40120;
  wire  T_40121;
  wire  T_40122;
  wire  T_40123;
  wire  T_40139;
  wire  T_40140;
  wire  T_40141;
  wire  T_40142;
  wire  T_40143;
  wire  T_40158;
  wire  T_40159;
  wire  T_40160;
  wire  T_40161;
  wire  T_40162;
  wire  T_40163;
  wire  T_40178;
  wire  T_40179;
  wire  T_40180;
  wire  T_40181;
  wire  T_40182;
  wire  T_40183;
  wire  T_40198;
  wire  T_40199;
  wire  T_40200;
  wire  T_40201;
  wire  T_40202;
  wire  T_40203;
  wire  T_40218;
  wire  T_40219;
  wire  T_40220;
  wire  T_40221;
  wire  T_40222;
  wire  T_40223;
  wire  T_40237;
  wire  T_40238;
  wire  T_40239;
  wire  T_40240;
  wire  T_40241;
  wire  T_40242;
  wire  T_40243;
  wire  T_40257;
  wire  T_40258;
  wire  T_40259;
  wire  T_40260;
  wire  T_40261;
  wire  T_40262;
  wire  T_40263;
  wire  T_40277;
  wire  T_40278;
  wire  T_40279;
  wire  T_40280;
  wire  T_40281;
  wire  T_40282;
  wire  T_40283;
  wire  T_40297;
  wire  T_40298;
  wire  T_40299;
  wire  T_40300;
  wire  T_40301;
  wire  T_40302;
  wire  T_40303;
  wire  T_40316;
  wire  T_40317;
  wire  T_40318;
  wire  T_40319;
  wire  T_40320;
  wire  T_40321;
  wire  T_40322;
  wire  T_40323;
  wire  T_40336;
  wire  T_40337;
  wire  T_40338;
  wire  T_40339;
  wire  T_40340;
  wire  T_40341;
  wire  T_40342;
  wire  T_40343;
  wire  T_40356;
  wire  T_40357;
  wire  T_40358;
  wire  T_40359;
  wire  T_40360;
  wire  T_40361;
  wire  T_40362;
  wire  T_40363;
  wire  T_40376;
  wire  T_40377;
  wire  T_40378;
  wire  T_40379;
  wire  T_40380;
  wire  T_40381;
  wire  T_40382;
  wire  T_40383;
  wire  T_40395;
  wire  T_40396;
  wire  T_40397;
  wire  T_40398;
  wire  T_40399;
  wire  T_40400;
  wire  T_40401;
  wire  T_40402;
  wire  T_40403;
  wire  T_40415;
  wire  T_40416;
  wire  T_40417;
  wire  T_40418;
  wire  T_40419;
  wire  T_40420;
  wire  T_40421;
  wire  T_40422;
  wire  T_40423;
  wire  T_40435;
  wire  T_40436;
  wire  T_40437;
  wire  T_40438;
  wire  T_40439;
  wire  T_40440;
  wire  T_40441;
  wire  T_40442;
  wire  T_40443;
  wire  T_40455;
  wire  T_40456;
  wire  T_40457;
  wire  T_40458;
  wire  T_40459;
  wire  T_40460;
  wire  T_40461;
  wire  T_40462;
  wire  T_40463;
  wire  T_40474;
  wire  T_40475;
  wire  T_40476;
  wire  T_40477;
  wire  T_40478;
  wire  T_40479;
  wire  T_40480;
  wire  T_40481;
  wire  T_40482;
  wire  T_40483;
  wire  T_40494;
  wire  T_40495;
  wire  T_40496;
  wire  T_40497;
  wire  T_40498;
  wire  T_40499;
  wire  T_40500;
  wire  T_40501;
  wire  T_40502;
  wire  T_40503;
  wire  T_40514;
  wire  T_40515;
  wire  T_40516;
  wire  T_40517;
  wire  T_40518;
  wire  T_40519;
  wire  T_40520;
  wire  T_40521;
  wire  T_40522;
  wire  T_40523;
  wire  T_40534;
  wire  T_40535;
  wire  T_40536;
  wire  T_40537;
  wire  T_40538;
  wire  T_40539;
  wire  T_40540;
  wire  T_40541;
  wire  T_40542;
  wire  T_40543;
  wire  T_40553;
  wire  T_40554;
  wire  T_40555;
  wire  T_40556;
  wire  T_40557;
  wire  T_40558;
  wire  T_40559;
  wire  T_40560;
  wire  T_40561;
  wire  T_40562;
  wire  T_40563;
  wire  T_40573;
  wire  T_40574;
  wire  T_40575;
  wire  T_40576;
  wire  T_40577;
  wire  T_40578;
  wire  T_40579;
  wire  T_40580;
  wire  T_40581;
  wire  T_40582;
  wire  T_40583;
  wire  T_40593;
  wire  T_40594;
  wire  T_40595;
  wire  T_40596;
  wire  T_40597;
  wire  T_40598;
  wire  T_40599;
  wire  T_40600;
  wire  T_40601;
  wire  T_40602;
  wire  T_40603;
  wire  T_40613;
  wire  T_40614;
  wire  T_40615;
  wire  T_40616;
  wire  T_40617;
  wire  T_40618;
  wire  T_40619;
  wire  T_40620;
  wire  T_40621;
  wire  T_40622;
  wire  T_40623;
  wire  T_40632;
  wire  T_40633;
  wire  T_40634;
  wire  T_40635;
  wire  T_40636;
  wire  T_40637;
  wire  T_40638;
  wire  T_40639;
  wire  T_40640;
  wire  T_40641;
  wire  T_40642;
  wire  T_40643;
  wire  T_40652;
  wire  T_40653;
  wire  T_40654;
  wire  T_40655;
  wire  T_40656;
  wire  T_40657;
  wire  T_40658;
  wire  T_40659;
  wire  T_40660;
  wire  T_40661;
  wire  T_40662;
  wire  T_40663;
  wire  T_40672;
  wire  T_40673;
  wire  T_40674;
  wire  T_40675;
  wire  T_40676;
  wire  T_40677;
  wire  T_40678;
  wire  T_40679;
  wire  T_40680;
  wire  T_40681;
  wire  T_40682;
  wire  T_40683;
  wire  T_40692;
  wire  T_40693;
  wire  T_40694;
  wire  T_40695;
  wire  T_40696;
  wire  T_40697;
  wire  T_40698;
  wire  T_40699;
  wire  T_40700;
  wire  T_40701;
  wire  T_40702;
  wire  T_40703;
  wire  T_40711;
  wire  T_40712;
  wire  T_40713;
  wire  T_40714;
  wire  T_40715;
  wire  T_40716;
  wire  T_40717;
  wire  T_40718;
  wire  T_40719;
  wire  T_40720;
  wire  T_40721;
  wire  T_40722;
  wire  T_40723;
  wire  T_40731;
  wire  T_40732;
  wire  T_40733;
  wire  T_40734;
  wire  T_40735;
  wire  T_40736;
  wire  T_40737;
  wire  T_40738;
  wire  T_40739;
  wire  T_40740;
  wire  T_40741;
  wire  T_40742;
  wire  T_40743;
  wire  T_40751;
  wire  T_40752;
  wire  T_40753;
  wire  T_40754;
  wire  T_40755;
  wire  T_40756;
  wire  T_40757;
  wire  T_40758;
  wire  T_40759;
  wire  T_40760;
  wire  T_40761;
  wire  T_40762;
  wire  T_40763;
  wire  T_40771;
  wire  T_40772;
  wire  T_40773;
  wire  T_40774;
  wire  T_40775;
  wire  T_40776;
  wire  T_40777;
  wire  T_40778;
  wire  T_40779;
  wire  T_40780;
  wire  T_40781;
  wire  T_40782;
  wire  T_40783;
  wire  T_40790;
  wire  T_40791;
  wire  T_40792;
  wire  T_40793;
  wire  T_40794;
  wire  T_40795;
  wire  T_40796;
  wire  T_40797;
  wire  T_40798;
  wire  T_40799;
  wire  T_40800;
  wire  T_40801;
  wire  T_40802;
  wire  T_40803;
  wire  T_40810;
  wire  T_40811;
  wire  T_40812;
  wire  T_40813;
  wire  T_40814;
  wire  T_40815;
  wire  T_40816;
  wire  T_40817;
  wire  T_40818;
  wire  T_40819;
  wire  T_40820;
  wire  T_40821;
  wire  T_40822;
  wire  T_40823;
  wire  T_40830;
  wire  T_40831;
  wire  T_40832;
  wire  T_40833;
  wire  T_40834;
  wire  T_40835;
  wire  T_40836;
  wire  T_40837;
  wire  T_40838;
  wire  T_40839;
  wire  T_40840;
  wire  T_40841;
  wire  T_40842;
  wire  T_40843;
  wire  T_40850;
  wire  T_40851;
  wire  T_40852;
  wire  T_40853;
  wire  T_40854;
  wire  T_40855;
  wire  T_40856;
  wire  T_40857;
  wire  T_40858;
  wire  T_40859;
  wire  T_40860;
  wire  T_40861;
  wire  T_40862;
  wire  T_40863;
  wire  T_40869;
  wire  T_40870;
  wire  T_40871;
  wire  T_40872;
  wire  T_40873;
  wire  T_40874;
  wire  T_40875;
  wire  T_40876;
  wire  T_40877;
  wire  T_40878;
  wire  T_40879;
  wire  T_40880;
  wire  T_40881;
  wire  T_40882;
  wire  T_40883;
  wire  T_40889;
  wire  T_40890;
  wire  T_40891;
  wire  T_40892;
  wire  T_40893;
  wire  T_40894;
  wire  T_40895;
  wire  T_40896;
  wire  T_40897;
  wire  T_40898;
  wire  T_40899;
  wire  T_40900;
  wire  T_40901;
  wire  T_40902;
  wire  T_40903;
  wire  T_40909;
  wire  T_40910;
  wire  T_40911;
  wire  T_40912;
  wire  T_40913;
  wire  T_40914;
  wire  T_40915;
  wire  T_40916;
  wire  T_40917;
  wire  T_40918;
  wire  T_40919;
  wire  T_40920;
  wire  T_40921;
  wire  T_40922;
  wire  T_40923;
  wire  T_40929;
  wire  T_40930;
  wire  T_40931;
  wire  T_40932;
  wire  T_40933;
  wire  T_40934;
  wire  T_40935;
  wire  T_40936;
  wire  T_40937;
  wire  T_40938;
  wire  T_40939;
  wire  T_40940;
  wire  T_40941;
  wire  T_40942;
  wire  T_40943;
  wire  T_40948;
  wire  T_40949;
  wire  T_40950;
  wire  T_40951;
  wire  T_40952;
  wire  T_40953;
  wire  T_40954;
  wire  T_40955;
  wire  T_40956;
  wire  T_40957;
  wire  T_40958;
  wire  T_40959;
  wire  T_40960;
  wire  T_40961;
  wire  T_40962;
  wire  T_40963;
  wire  T_40968;
  wire  T_40969;
  wire  T_40970;
  wire  T_40971;
  wire  T_40972;
  wire  T_40973;
  wire  T_40974;
  wire  T_40975;
  wire  T_40976;
  wire  T_40977;
  wire  T_40978;
  wire  T_40979;
  wire  T_40980;
  wire  T_40981;
  wire  T_40982;
  wire  T_40983;
  wire  T_40988;
  wire  T_40989;
  wire  T_40990;
  wire  T_40991;
  wire  T_40992;
  wire  T_40993;
  wire  T_40994;
  wire  T_40995;
  wire  T_40996;
  wire  T_40997;
  wire  T_40998;
  wire  T_40999;
  wire  T_41000;
  wire  T_41001;
  wire  T_41002;
  wire  T_41003;
  wire  T_41008;
  wire  T_41009;
  wire  T_41010;
  wire  T_41011;
  wire  T_41012;
  wire  T_41013;
  wire  T_41014;
  wire  T_41015;
  wire  T_41016;
  wire  T_41017;
  wire  T_41018;
  wire  T_41019;
  wire  T_41020;
  wire  T_41021;
  wire  T_41022;
  wire  T_41023;
  wire  T_41027;
  wire  T_41028;
  wire  T_41029;
  wire  T_41030;
  wire  T_41031;
  wire  T_41032;
  wire  T_41033;
  wire  T_41034;
  wire  T_41035;
  wire  T_41036;
  wire  T_41037;
  wire  T_41038;
  wire  T_41039;
  wire  T_41040;
  wire  T_41041;
  wire  T_41042;
  wire  T_41043;
  wire  T_41047;
  wire  T_41048;
  wire  T_41049;
  wire  T_41050;
  wire  T_41051;
  wire  T_41052;
  wire  T_41053;
  wire  T_41054;
  wire  T_41055;
  wire  T_41056;
  wire  T_41057;
  wire  T_41058;
  wire  T_41059;
  wire  T_41060;
  wire  T_41061;
  wire  T_41062;
  wire  T_41063;
  wire  T_41067;
  wire  T_41068;
  wire  T_41069;
  wire  T_41070;
  wire  T_41071;
  wire  T_41072;
  wire  T_41073;
  wire  T_41074;
  wire  T_41075;
  wire  T_41076;
  wire  T_41077;
  wire  T_41078;
  wire  T_41079;
  wire  T_41080;
  wire  T_41081;
  wire  T_41082;
  wire  T_41083;
  wire  T_41087;
  wire  T_41088;
  wire  T_41089;
  wire  T_41090;
  wire  T_41091;
  wire  T_41092;
  wire  T_41093;
  wire  T_41094;
  wire  T_41095;
  wire  T_41096;
  wire  T_41097;
  wire  T_41098;
  wire  T_41099;
  wire  T_41100;
  wire  T_41101;
  wire  T_41102;
  wire  T_41103;
  wire  T_41106;
  wire  T_41107;
  wire  T_41108;
  wire  T_41109;
  wire  T_41110;
  wire  T_41111;
  wire  T_41112;
  wire  T_41113;
  wire  T_41114;
  wire  T_41115;
  wire  T_41116;
  wire  T_41117;
  wire  T_41118;
  wire  T_41119;
  wire  T_41120;
  wire  T_41121;
  wire  T_41122;
  wire  T_41123;
  wire  T_41126;
  wire  T_41127;
  wire  T_41128;
  wire  T_41129;
  wire  T_41130;
  wire  T_41131;
  wire  T_41132;
  wire  T_41133;
  wire  T_41134;
  wire  T_41135;
  wire  T_41136;
  wire  T_41137;
  wire  T_41138;
  wire  T_41139;
  wire  T_41140;
  wire  T_41141;
  wire  T_41142;
  wire  T_41143;
  wire  T_41146;
  wire  T_41147;
  wire  T_41148;
  wire  T_41149;
  wire  T_41150;
  wire  T_41151;
  wire  T_41152;
  wire  T_41153;
  wire  T_41154;
  wire  T_41155;
  wire  T_41156;
  wire  T_41157;
  wire  T_41158;
  wire  T_41159;
  wire  T_41160;
  wire  T_41161;
  wire  T_41162;
  wire  T_41163;
  wire  T_41166;
  wire  T_41167;
  wire  T_41168;
  wire  T_41169;
  wire  T_41170;
  wire  T_41171;
  wire  T_41172;
  wire  T_41173;
  wire  T_41174;
  wire  T_41175;
  wire  T_41176;
  wire  T_41177;
  wire  T_41178;
  wire  T_41179;
  wire  T_41180;
  wire  T_41181;
  wire  T_41182;
  wire  T_41183;
  wire  T_41185;
  wire  T_41186;
  wire  T_41187;
  wire  T_41188;
  wire  T_41189;
  wire  T_41190;
  wire  T_41191;
  wire  T_41192;
  wire  T_41193;
  wire  T_41194;
  wire  T_41195;
  wire  T_41196;
  wire  T_41197;
  wire  T_41198;
  wire  T_41199;
  wire  T_41200;
  wire  T_41201;
  wire  T_41202;
  wire  T_41203;
  wire  T_41205;
  wire  T_41206;
  wire  T_41207;
  wire  T_41208;
  wire  T_41209;
  wire  T_41210;
  wire  T_41211;
  wire  T_41212;
  wire  T_41213;
  wire  T_41214;
  wire  T_41215;
  wire  T_41216;
  wire  T_41217;
  wire  T_41218;
  wire  T_41219;
  wire  T_41220;
  wire  T_41221;
  wire  T_41222;
  wire  T_41223;
  wire  T_41225;
  wire  T_41226;
  wire  T_41227;
  wire  T_41228;
  wire  T_41229;
  wire  T_41230;
  wire  T_41231;
  wire  T_41232;
  wire  T_41233;
  wire  T_41234;
  wire  T_41235;
  wire  T_41236;
  wire  T_41237;
  wire  T_41238;
  wire  T_41239;
  wire  T_41240;
  wire  T_41241;
  wire  T_41242;
  wire  T_41243;
  wire  T_41245;
  wire  T_41246;
  wire  T_41247;
  wire  T_41248;
  wire  T_41249;
  wire  T_41250;
  wire  T_41251;
  wire  T_41252;
  wire  T_41253;
  wire  T_41254;
  wire  T_41255;
  wire  T_41256;
  wire  T_41257;
  wire  T_41258;
  wire  T_41259;
  wire  T_41260;
  wire  T_41261;
  wire  T_41262;
  wire  T_41263;
  wire  T_41337;
  wire  T_41338;
  wire  T_41339;
  wire  T_41340;
  wire  T_41341;
  wire  T_41342;
  wire  T_41343;
  wire  T_41344;
  wire  T_41345;
  wire  T_41346;
  wire  T_41347;
  wire  T_41348;
  wire  T_41349;
  wire  T_41350;
  wire  T_41351;
  wire  T_41352;
  wire  T_41353;
  wire  T_41354;
  wire  T_41355;
  wire  T_41356;
  wire  T_41357;
  wire  T_41358;
  wire  T_41359;
  wire  T_41360;
  wire  T_41361;
  wire  T_41362;
  wire  T_41363;
  wire  T_41364;
  wire  T_41365;
  wire  T_41366;
  wire  T_41367;
  wire  T_41369;
  wire  T_41370;
  wire  T_41371;
  wire  T_41372;
  wire  T_41373;
  wire  T_41374;
  wire  T_41375;
  wire  T_41376;
  wire  T_41377;
  wire  T_41378;
  wire  T_41379;
  wire  T_41380;
  wire  T_41381;
  wire  T_41382;
  wire  T_41383;
  wire  T_41384;
  wire  T_41385;
  wire  T_41386;
  wire  T_41387;
  wire  T_41388;
  wire  T_41389;
  wire  T_41390;
  wire  T_41391;
  wire  T_41392;
  wire  T_41393;
  wire  T_41394;
  wire  T_41395;
  wire  T_41396;
  wire  T_41397;
  wire  T_41398;
  wire  T_41399;
  wire  T_41401;
  wire  T_41402;
  wire  T_41403;
  wire  T_41404;
  wire  T_41405;
  wire  T_41406;
  wire  T_41407;
  wire  T_41408;
  wire  T_41409;
  wire  T_41410;
  wire  T_41411;
  wire  T_41412;
  wire  T_41413;
  wire  T_41414;
  wire  T_41415;
  wire  T_41416;
  wire  T_41417;
  wire  T_41418;
  wire  T_41419;
  wire  T_41420;
  wire  T_41421;
  wire  T_41422;
  wire  T_41423;
  wire  T_41424;
  wire  T_41425;
  wire  T_41426;
  wire  T_41427;
  wire  T_41428;
  wire  T_41429;
  wire  T_41430;
  wire  T_41431;
  wire  T_41433;
  wire  T_41434;
  wire  T_41435;
  wire  T_41436;
  wire  T_41437;
  wire  T_41438;
  wire  T_41439;
  wire  T_41440;
  wire  T_41441;
  wire  T_41442;
  wire  T_41443;
  wire  T_41444;
  wire  T_41445;
  wire  T_41446;
  wire  T_41447;
  wire  T_41448;
  wire  T_41449;
  wire  T_41450;
  wire  T_41451;
  wire  T_41452;
  wire  T_41453;
  wire  T_41454;
  wire  T_41455;
  wire  T_41456;
  wire  T_41457;
  wire  T_41458;
  wire  T_41459;
  wire  T_41460;
  wire  T_41461;
  wire  T_41462;
  wire  T_41463;
  wire  T_41495;
  wire  T_41527;
  wire  T_41559;
  wire  T_41591;
  wire  T_41622;
  wire  T_41623;
  wire  T_41654;
  wire  T_41655;
  wire  T_41686;
  wire  T_41687;
  wire  T_41718;
  wire  T_41719;
  wire  T_41749;
  wire  T_41750;
  wire  T_41751;
  wire  T_41781;
  wire  T_41782;
  wire  T_41783;
  wire  T_41813;
  wire  T_41814;
  wire  T_41815;
  wire  T_41845;
  wire  T_41846;
  wire  T_41847;
  wire  T_41876;
  wire  T_41877;
  wire  T_41878;
  wire  T_41879;
  wire  T_41908;
  wire  T_41909;
  wire  T_41910;
  wire  T_41911;
  wire  T_41940;
  wire  T_41941;
  wire  T_41942;
  wire  T_41943;
  wire  T_41972;
  wire  T_41973;
  wire  T_41974;
  wire  T_41975;
  wire  T_42003;
  wire  T_42004;
  wire  T_42005;
  wire  T_42006;
  wire  T_42007;
  wire  T_42035;
  wire  T_42036;
  wire  T_42037;
  wire  T_42038;
  wire  T_42039;
  wire  T_42067;
  wire  T_42068;
  wire  T_42069;
  wire  T_42070;
  wire  T_42071;
  wire  T_42099;
  wire  T_42100;
  wire  T_42101;
  wire  T_42102;
  wire  T_42103;
  wire  T_42130;
  wire  T_42131;
  wire  T_42132;
  wire  T_42133;
  wire  T_42134;
  wire  T_42135;
  wire  T_42162;
  wire  T_42163;
  wire  T_42164;
  wire  T_42165;
  wire  T_42166;
  wire  T_42167;
  wire  T_42194;
  wire  T_42195;
  wire  T_42196;
  wire  T_42197;
  wire  T_42198;
  wire  T_42199;
  wire  T_42226;
  wire  T_42227;
  wire  T_42228;
  wire  T_42229;
  wire  T_42230;
  wire  T_42231;
  wire  T_42257;
  wire  T_42258;
  wire  T_42259;
  wire  T_42260;
  wire  T_42261;
  wire  T_42262;
  wire  T_42263;
  wire  T_42289;
  wire  T_42290;
  wire  T_42291;
  wire  T_42292;
  wire  T_42293;
  wire  T_42294;
  wire  T_42295;
  wire  T_42321;
  wire  T_42322;
  wire  T_42323;
  wire  T_42324;
  wire  T_42325;
  wire  T_42326;
  wire  T_42327;
  wire  T_42353;
  wire  T_42354;
  wire  T_42355;
  wire  T_42356;
  wire  T_42357;
  wire  T_42358;
  wire  T_42359;
  wire  T_42384;
  wire  T_42385;
  wire  T_42386;
  wire  T_42387;
  wire  T_42388;
  wire  T_42389;
  wire  T_42390;
  wire  T_42391;
  wire  T_42416;
  wire  T_42417;
  wire  T_42418;
  wire  T_42419;
  wire  T_42420;
  wire  T_42421;
  wire  T_42422;
  wire  T_42423;
  wire  T_42448;
  wire  T_42449;
  wire  T_42450;
  wire  T_42451;
  wire  T_42452;
  wire  T_42453;
  wire  T_42454;
  wire  T_42455;
  wire  T_42480;
  wire  T_42481;
  wire  T_42482;
  wire  T_42483;
  wire  T_42484;
  wire  T_42485;
  wire  T_42486;
  wire  T_42487;
  wire  T_42511;
  wire  T_42512;
  wire  T_42513;
  wire  T_42514;
  wire  T_42515;
  wire  T_42516;
  wire  T_42517;
  wire  T_42518;
  wire  T_42519;
  wire  T_42543;
  wire  T_42544;
  wire  T_42545;
  wire  T_42546;
  wire  T_42547;
  wire  T_42548;
  wire  T_42549;
  wire  T_42550;
  wire  T_42551;
  wire  T_42575;
  wire  T_42576;
  wire  T_42577;
  wire  T_42578;
  wire  T_42579;
  wire  T_42580;
  wire  T_42581;
  wire  T_42582;
  wire  T_42583;
  wire  T_42607;
  wire  T_42608;
  wire  T_42609;
  wire  T_42610;
  wire  T_42611;
  wire  T_42612;
  wire  T_42613;
  wire  T_42614;
  wire  T_42615;
  wire  T_42638;
  wire  T_42639;
  wire  T_42640;
  wire  T_42641;
  wire  T_42642;
  wire  T_42643;
  wire  T_42644;
  wire  T_42645;
  wire  T_42646;
  wire  T_42647;
  wire  T_42670;
  wire  T_42671;
  wire  T_42672;
  wire  T_42673;
  wire  T_42674;
  wire  T_42675;
  wire  T_42676;
  wire  T_42677;
  wire  T_42678;
  wire  T_42679;
  wire  T_42702;
  wire  T_42703;
  wire  T_42704;
  wire  T_42705;
  wire  T_42706;
  wire  T_42707;
  wire  T_42708;
  wire  T_42709;
  wire  T_42710;
  wire  T_42711;
  wire  T_42734;
  wire  T_42735;
  wire  T_42736;
  wire  T_42737;
  wire  T_42738;
  wire  T_42739;
  wire  T_42740;
  wire  T_42741;
  wire  T_42742;
  wire  T_42743;
  wire  T_42765;
  wire  T_42766;
  wire  T_42767;
  wire  T_42768;
  wire  T_42769;
  wire  T_42770;
  wire  T_42771;
  wire  T_42772;
  wire  T_42773;
  wire  T_42774;
  wire  T_42775;
  wire  T_42797;
  wire  T_42798;
  wire  T_42799;
  wire  T_42800;
  wire  T_42801;
  wire  T_42802;
  wire  T_42803;
  wire  T_42804;
  wire  T_42805;
  wire  T_42806;
  wire  T_42807;
  wire  T_42829;
  wire  T_42830;
  wire  T_42831;
  wire  T_42832;
  wire  T_42833;
  wire  T_42834;
  wire  T_42835;
  wire  T_42836;
  wire  T_42837;
  wire  T_42838;
  wire  T_42839;
  wire  T_42861;
  wire  T_42862;
  wire  T_42863;
  wire  T_42864;
  wire  T_42865;
  wire  T_42866;
  wire  T_42867;
  wire  T_42868;
  wire  T_42869;
  wire  T_42870;
  wire  T_42871;
  wire  T_42892;
  wire  T_42893;
  wire  T_42894;
  wire  T_42895;
  wire  T_42896;
  wire  T_42897;
  wire  T_42898;
  wire  T_42899;
  wire  T_42900;
  wire  T_42901;
  wire  T_42902;
  wire  T_42903;
  wire  T_42924;
  wire  T_42925;
  wire  T_42926;
  wire  T_42927;
  wire  T_42928;
  wire  T_42929;
  wire  T_42930;
  wire  T_42931;
  wire  T_42932;
  wire  T_42933;
  wire  T_42934;
  wire  T_42935;
  wire  T_42956;
  wire  T_42957;
  wire  T_42958;
  wire  T_42959;
  wire  T_42960;
  wire  T_42961;
  wire  T_42962;
  wire  T_42963;
  wire  T_42964;
  wire  T_42965;
  wire  T_42966;
  wire  T_42967;
  wire  T_42988;
  wire  T_42989;
  wire  T_42990;
  wire  T_42991;
  wire  T_42992;
  wire  T_42993;
  wire  T_42994;
  wire  T_42995;
  wire  T_42996;
  wire  T_42997;
  wire  T_42998;
  wire  T_42999;
  wire  T_43019;
  wire  T_43020;
  wire  T_43021;
  wire  T_43022;
  wire  T_43023;
  wire  T_43024;
  wire  T_43025;
  wire  T_43026;
  wire  T_43027;
  wire  T_43028;
  wire  T_43029;
  wire  T_43030;
  wire  T_43031;
  wire  T_43051;
  wire  T_43052;
  wire  T_43053;
  wire  T_43054;
  wire  T_43055;
  wire  T_43056;
  wire  T_43057;
  wire  T_43058;
  wire  T_43059;
  wire  T_43060;
  wire  T_43061;
  wire  T_43062;
  wire  T_43063;
  wire  T_43083;
  wire  T_43084;
  wire  T_43085;
  wire  T_43086;
  wire  T_43087;
  wire  T_43088;
  wire  T_43089;
  wire  T_43090;
  wire  T_43091;
  wire  T_43092;
  wire  T_43093;
  wire  T_43094;
  wire  T_43095;
  wire  T_43115;
  wire  T_43116;
  wire  T_43117;
  wire  T_43118;
  wire  T_43119;
  wire  T_43120;
  wire  T_43121;
  wire  T_43122;
  wire  T_43123;
  wire  T_43124;
  wire  T_43125;
  wire  T_43126;
  wire  T_43127;
  wire  T_43146;
  wire  T_43147;
  wire  T_43148;
  wire  T_43149;
  wire  T_43150;
  wire  T_43151;
  wire  T_43152;
  wire  T_43153;
  wire  T_43154;
  wire  T_43155;
  wire  T_43156;
  wire  T_43157;
  wire  T_43158;
  wire  T_43159;
  wire  T_43178;
  wire  T_43179;
  wire  T_43180;
  wire  T_43181;
  wire  T_43182;
  wire  T_43183;
  wire  T_43184;
  wire  T_43185;
  wire  T_43186;
  wire  T_43187;
  wire  T_43188;
  wire  T_43189;
  wire  T_43190;
  wire  T_43191;
  wire  T_43210;
  wire  T_43211;
  wire  T_43212;
  wire  T_43213;
  wire  T_43214;
  wire  T_43215;
  wire  T_43216;
  wire  T_43217;
  wire  T_43218;
  wire  T_43219;
  wire  T_43220;
  wire  T_43221;
  wire  T_43222;
  wire  T_43223;
  wire  T_43242;
  wire  T_43243;
  wire  T_43244;
  wire  T_43245;
  wire  T_43246;
  wire  T_43247;
  wire  T_43248;
  wire  T_43249;
  wire  T_43250;
  wire  T_43251;
  wire  T_43252;
  wire  T_43253;
  wire  T_43254;
  wire  T_43255;
  wire  T_43273;
  wire  T_43274;
  wire  T_43275;
  wire  T_43276;
  wire  T_43277;
  wire  T_43278;
  wire  T_43279;
  wire  T_43280;
  wire  T_43281;
  wire  T_43282;
  wire  T_43283;
  wire  T_43284;
  wire  T_43285;
  wire  T_43286;
  wire  T_43287;
  wire  T_43305;
  wire  T_43306;
  wire  T_43307;
  wire  T_43308;
  wire  T_43309;
  wire  T_43310;
  wire  T_43311;
  wire  T_43312;
  wire  T_43313;
  wire  T_43314;
  wire  T_43315;
  wire  T_43316;
  wire  T_43317;
  wire  T_43318;
  wire  T_43319;
  wire  T_43337;
  wire  T_43338;
  wire  T_43339;
  wire  T_43340;
  wire  T_43341;
  wire  T_43342;
  wire  T_43343;
  wire  T_43344;
  wire  T_43345;
  wire  T_43346;
  wire  T_43347;
  wire  T_43348;
  wire  T_43349;
  wire  T_43350;
  wire  T_43351;
  wire  T_43369;
  wire  T_43370;
  wire  T_43371;
  wire  T_43372;
  wire  T_43373;
  wire  T_43374;
  wire  T_43375;
  wire  T_43376;
  wire  T_43377;
  wire  T_43378;
  wire  T_43379;
  wire  T_43380;
  wire  T_43381;
  wire  T_43382;
  wire  T_43383;
  wire  T_43400;
  wire  T_43401;
  wire  T_43402;
  wire  T_43403;
  wire  T_43404;
  wire  T_43405;
  wire  T_43406;
  wire  T_43407;
  wire  T_43408;
  wire  T_43409;
  wire  T_43410;
  wire  T_43411;
  wire  T_43412;
  wire  T_43413;
  wire  T_43414;
  wire  T_43415;
  wire  T_43432;
  wire  T_43433;
  wire  T_43434;
  wire  T_43435;
  wire  T_43436;
  wire  T_43437;
  wire  T_43438;
  wire  T_43439;
  wire  T_43440;
  wire  T_43441;
  wire  T_43442;
  wire  T_43443;
  wire  T_43444;
  wire  T_43445;
  wire  T_43446;
  wire  T_43447;
  wire  T_43464;
  wire  T_43465;
  wire  T_43466;
  wire  T_43467;
  wire  T_43468;
  wire  T_43469;
  wire  T_43470;
  wire  T_43471;
  wire  T_43472;
  wire  T_43473;
  wire  T_43474;
  wire  T_43475;
  wire  T_43476;
  wire  T_43477;
  wire  T_43478;
  wire  T_43479;
  wire  T_43496;
  wire  T_43497;
  wire  T_43498;
  wire  T_43499;
  wire  T_43500;
  wire  T_43501;
  wire  T_43502;
  wire  T_43503;
  wire  T_43504;
  wire  T_43505;
  wire  T_43506;
  wire  T_43507;
  wire  T_43508;
  wire  T_43509;
  wire  T_43510;
  wire  T_43511;
  wire  T_43527;
  wire  T_43528;
  wire  T_43529;
  wire  T_43530;
  wire  T_43531;
  wire  T_43532;
  wire  T_43533;
  wire  T_43534;
  wire  T_43535;
  wire  T_43536;
  wire  T_43537;
  wire  T_43538;
  wire  T_43539;
  wire  T_43540;
  wire  T_43541;
  wire  T_43542;
  wire  T_43543;
  wire  T_43559;
  wire  T_43560;
  wire  T_43561;
  wire  T_43562;
  wire  T_43563;
  wire  T_43564;
  wire  T_43565;
  wire  T_43566;
  wire  T_43567;
  wire  T_43568;
  wire  T_43569;
  wire  T_43570;
  wire  T_43571;
  wire  T_43572;
  wire  T_43573;
  wire  T_43574;
  wire  T_43575;
  wire  T_43591;
  wire  T_43592;
  wire  T_43593;
  wire  T_43594;
  wire  T_43595;
  wire  T_43596;
  wire  T_43597;
  wire  T_43598;
  wire  T_43599;
  wire  T_43600;
  wire  T_43601;
  wire  T_43602;
  wire  T_43603;
  wire  T_43604;
  wire  T_43605;
  wire  T_43606;
  wire  T_43607;
  wire  T_43623;
  wire  T_43624;
  wire  T_43625;
  wire  T_43626;
  wire  T_43627;
  wire  T_43628;
  wire  T_43629;
  wire  T_43630;
  wire  T_43631;
  wire  T_43632;
  wire  T_43633;
  wire  T_43634;
  wire  T_43635;
  wire  T_43636;
  wire  T_43637;
  wire  T_43638;
  wire  T_43639;
  wire  T_43654;
  wire  T_43655;
  wire  T_43656;
  wire  T_43657;
  wire  T_43658;
  wire  T_43659;
  wire  T_43660;
  wire  T_43661;
  wire  T_43662;
  wire  T_43663;
  wire  T_43664;
  wire  T_43665;
  wire  T_43666;
  wire  T_43667;
  wire  T_43668;
  wire  T_43669;
  wire  T_43670;
  wire  T_43671;
  wire  T_43686;
  wire  T_43687;
  wire  T_43688;
  wire  T_43689;
  wire  T_43690;
  wire  T_43691;
  wire  T_43692;
  wire  T_43693;
  wire  T_43694;
  wire  T_43695;
  wire  T_43696;
  wire  T_43697;
  wire  T_43698;
  wire  T_43699;
  wire  T_43700;
  wire  T_43701;
  wire  T_43702;
  wire  T_43703;
  wire  T_43718;
  wire  T_43719;
  wire  T_43720;
  wire  T_43721;
  wire  T_43722;
  wire  T_43723;
  wire  T_43724;
  wire  T_43725;
  wire  T_43726;
  wire  T_43727;
  wire  T_43728;
  wire  T_43729;
  wire  T_43730;
  wire  T_43731;
  wire  T_43732;
  wire  T_43733;
  wire  T_43734;
  wire  T_43735;
  wire  T_43750;
  wire  T_43751;
  wire  T_43752;
  wire  T_43753;
  wire  T_43754;
  wire  T_43755;
  wire  T_43756;
  wire  T_43757;
  wire  T_43758;
  wire  T_43759;
  wire  T_43760;
  wire  T_43761;
  wire  T_43762;
  wire  T_43763;
  wire  T_43764;
  wire  T_43765;
  wire  T_43766;
  wire  T_43767;
  wire  T_43781;
  wire  T_43782;
  wire  T_43783;
  wire  T_43784;
  wire  T_43785;
  wire  T_43786;
  wire  T_43787;
  wire  T_43788;
  wire  T_43789;
  wire  T_43790;
  wire  T_43791;
  wire  T_43792;
  wire  T_43793;
  wire  T_43794;
  wire  T_43795;
  wire  T_43796;
  wire  T_43797;
  wire  T_43798;
  wire  T_43799;
  wire  T_43813;
  wire  T_43814;
  wire  T_43815;
  wire  T_43816;
  wire  T_43817;
  wire  T_43818;
  wire  T_43819;
  wire  T_43820;
  wire  T_43821;
  wire  T_43822;
  wire  T_43823;
  wire  T_43824;
  wire  T_43825;
  wire  T_43826;
  wire  T_43827;
  wire  T_43828;
  wire  T_43829;
  wire  T_43830;
  wire  T_43831;
  wire  T_43845;
  wire  T_43846;
  wire  T_43847;
  wire  T_43848;
  wire  T_43849;
  wire  T_43850;
  wire  T_43851;
  wire  T_43852;
  wire  T_43853;
  wire  T_43854;
  wire  T_43855;
  wire  T_43856;
  wire  T_43857;
  wire  T_43858;
  wire  T_43859;
  wire  T_43860;
  wire  T_43861;
  wire  T_43862;
  wire  T_43863;
  wire  T_43877;
  wire  T_43878;
  wire  T_43879;
  wire  T_43880;
  wire  T_43881;
  wire  T_43882;
  wire  T_43883;
  wire  T_43884;
  wire  T_43885;
  wire  T_43886;
  wire  T_43887;
  wire  T_43888;
  wire  T_43889;
  wire  T_43890;
  wire  T_43891;
  wire  T_43892;
  wire  T_43893;
  wire  T_43894;
  wire  T_43895;
  wire  T_43908;
  wire  T_43909;
  wire  T_43910;
  wire  T_43911;
  wire  T_43912;
  wire  T_43913;
  wire  T_43914;
  wire  T_43915;
  wire  T_43916;
  wire  T_43917;
  wire  T_43918;
  wire  T_43919;
  wire  T_43920;
  wire  T_43921;
  wire  T_43922;
  wire  T_43923;
  wire  T_43924;
  wire  T_43925;
  wire  T_43926;
  wire  T_43927;
  wire  T_43940;
  wire  T_43941;
  wire  T_43942;
  wire  T_43943;
  wire  T_43944;
  wire  T_43945;
  wire  T_43946;
  wire  T_43947;
  wire  T_43948;
  wire  T_43949;
  wire  T_43950;
  wire  T_43951;
  wire  T_43952;
  wire  T_43953;
  wire  T_43954;
  wire  T_43955;
  wire  T_43956;
  wire  T_43957;
  wire  T_43958;
  wire  T_43959;
  wire  T_43972;
  wire  T_43973;
  wire  T_43974;
  wire  T_43975;
  wire  T_43976;
  wire  T_43977;
  wire  T_43978;
  wire  T_43979;
  wire  T_43980;
  wire  T_43981;
  wire  T_43982;
  wire  T_43983;
  wire  T_43984;
  wire  T_43985;
  wire  T_43986;
  wire  T_43987;
  wire  T_43988;
  wire  T_43989;
  wire  T_43990;
  wire  T_43991;
  wire  T_44004;
  wire  T_44005;
  wire  T_44006;
  wire  T_44007;
  wire  T_44008;
  wire  T_44009;
  wire  T_44010;
  wire  T_44011;
  wire  T_44012;
  wire  T_44013;
  wire  T_44014;
  wire  T_44015;
  wire  T_44016;
  wire  T_44017;
  wire  T_44018;
  wire  T_44019;
  wire  T_44020;
  wire  T_44021;
  wire  T_44022;
  wire  T_44023;
  wire  T_44035;
  wire  T_44036;
  wire  T_44037;
  wire  T_44038;
  wire  T_44039;
  wire  T_44040;
  wire  T_44041;
  wire  T_44042;
  wire  T_44043;
  wire  T_44044;
  wire  T_44045;
  wire  T_44046;
  wire  T_44047;
  wire  T_44048;
  wire  T_44049;
  wire  T_44050;
  wire  T_44051;
  wire  T_44052;
  wire  T_44053;
  wire  T_44054;
  wire  T_44055;
  wire  T_44067;
  wire  T_44068;
  wire  T_44069;
  wire  T_44070;
  wire  T_44071;
  wire  T_44072;
  wire  T_44073;
  wire  T_44074;
  wire  T_44075;
  wire  T_44076;
  wire  T_44077;
  wire  T_44078;
  wire  T_44079;
  wire  T_44080;
  wire  T_44081;
  wire  T_44082;
  wire  T_44083;
  wire  T_44084;
  wire  T_44085;
  wire  T_44086;
  wire  T_44087;
  wire  T_44099;
  wire  T_44100;
  wire  T_44101;
  wire  T_44102;
  wire  T_44103;
  wire  T_44104;
  wire  T_44105;
  wire  T_44106;
  wire  T_44107;
  wire  T_44108;
  wire  T_44109;
  wire  T_44110;
  wire  T_44111;
  wire  T_44112;
  wire  T_44113;
  wire  T_44114;
  wire  T_44115;
  wire  T_44116;
  wire  T_44117;
  wire  T_44118;
  wire  T_44119;
  wire  T_44131;
  wire  T_44132;
  wire  T_44133;
  wire  T_44134;
  wire  T_44135;
  wire  T_44136;
  wire  T_44137;
  wire  T_44138;
  wire  T_44139;
  wire  T_44140;
  wire  T_44141;
  wire  T_44142;
  wire  T_44143;
  wire  T_44144;
  wire  T_44145;
  wire  T_44146;
  wire  T_44147;
  wire  T_44148;
  wire  T_44149;
  wire  T_44150;
  wire  T_44151;
  wire  T_44162;
  wire  T_44163;
  wire  T_44164;
  wire  T_44165;
  wire  T_44166;
  wire  T_44167;
  wire  T_44168;
  wire  T_44169;
  wire  T_44170;
  wire  T_44171;
  wire  T_44172;
  wire  T_44173;
  wire  T_44174;
  wire  T_44175;
  wire  T_44176;
  wire  T_44177;
  wire  T_44178;
  wire  T_44179;
  wire  T_44180;
  wire  T_44181;
  wire  T_44182;
  wire  T_44183;
  wire  T_44194;
  wire  T_44195;
  wire  T_44196;
  wire  T_44197;
  wire  T_44198;
  wire  T_44199;
  wire  T_44200;
  wire  T_44201;
  wire  T_44202;
  wire  T_44203;
  wire  T_44204;
  wire  T_44205;
  wire  T_44206;
  wire  T_44207;
  wire  T_44208;
  wire  T_44209;
  wire  T_44210;
  wire  T_44211;
  wire  T_44212;
  wire  T_44213;
  wire  T_44214;
  wire  T_44215;
  wire  T_44226;
  wire  T_44227;
  wire  T_44228;
  wire  T_44229;
  wire  T_44230;
  wire  T_44231;
  wire  T_44232;
  wire  T_44233;
  wire  T_44234;
  wire  T_44235;
  wire  T_44236;
  wire  T_44237;
  wire  T_44238;
  wire  T_44239;
  wire  T_44240;
  wire  T_44241;
  wire  T_44242;
  wire  T_44243;
  wire  T_44244;
  wire  T_44245;
  wire  T_44246;
  wire  T_44247;
  wire  T_44258;
  wire  T_44259;
  wire  T_44260;
  wire  T_44261;
  wire  T_44262;
  wire  T_44263;
  wire  T_44264;
  wire  T_44265;
  wire  T_44266;
  wire  T_44267;
  wire  T_44268;
  wire  T_44269;
  wire  T_44270;
  wire  T_44271;
  wire  T_44272;
  wire  T_44273;
  wire  T_44274;
  wire  T_44275;
  wire  T_44276;
  wire  T_44277;
  wire  T_44278;
  wire  T_44279;
  wire  T_44289;
  wire  T_44290;
  wire  T_44291;
  wire  T_44292;
  wire  T_44293;
  wire  T_44294;
  wire  T_44295;
  wire  T_44296;
  wire  T_44297;
  wire  T_44298;
  wire  T_44299;
  wire  T_44300;
  wire  T_44301;
  wire  T_44302;
  wire  T_44303;
  wire  T_44304;
  wire  T_44305;
  wire  T_44306;
  wire  T_44307;
  wire  T_44308;
  wire  T_44309;
  wire  T_44310;
  wire  T_44311;
  wire  T_44321;
  wire  T_44322;
  wire  T_44323;
  wire  T_44324;
  wire  T_44325;
  wire  T_44326;
  wire  T_44327;
  wire  T_44328;
  wire  T_44329;
  wire  T_44330;
  wire  T_44331;
  wire  T_44332;
  wire  T_44333;
  wire  T_44334;
  wire  T_44335;
  wire  T_44336;
  wire  T_44337;
  wire  T_44338;
  wire  T_44339;
  wire  T_44340;
  wire  T_44341;
  wire  T_44342;
  wire  T_44343;
  wire  T_44353;
  wire  T_44354;
  wire  T_44355;
  wire  T_44356;
  wire  T_44357;
  wire  T_44358;
  wire  T_44359;
  wire  T_44360;
  wire  T_44361;
  wire  T_44362;
  wire  T_44363;
  wire  T_44364;
  wire  T_44365;
  wire  T_44366;
  wire  T_44367;
  wire  T_44368;
  wire  T_44369;
  wire  T_44370;
  wire  T_44371;
  wire  T_44372;
  wire  T_44373;
  wire  T_44374;
  wire  T_44375;
  wire  T_44385;
  wire  T_44386;
  wire  T_44387;
  wire  T_44388;
  wire  T_44389;
  wire  T_44390;
  wire  T_44391;
  wire  T_44392;
  wire  T_44393;
  wire  T_44394;
  wire  T_44395;
  wire  T_44396;
  wire  T_44397;
  wire  T_44398;
  wire  T_44399;
  wire  T_44400;
  wire  T_44401;
  wire  T_44402;
  wire  T_44403;
  wire  T_44404;
  wire  T_44405;
  wire  T_44406;
  wire  T_44407;
  wire  T_44416;
  wire  T_44417;
  wire  T_44418;
  wire  T_44419;
  wire  T_44420;
  wire  T_44421;
  wire  T_44422;
  wire  T_44423;
  wire  T_44424;
  wire  T_44425;
  wire  T_44426;
  wire  T_44427;
  wire  T_44428;
  wire  T_44429;
  wire  T_44430;
  wire  T_44431;
  wire  T_44432;
  wire  T_44433;
  wire  T_44434;
  wire  T_44435;
  wire  T_44436;
  wire  T_44437;
  wire  T_44438;
  wire  T_44439;
  wire  T_44448;
  wire  T_44449;
  wire  T_44450;
  wire  T_44451;
  wire  T_44452;
  wire  T_44453;
  wire  T_44454;
  wire  T_44455;
  wire  T_44456;
  wire  T_44457;
  wire  T_44458;
  wire  T_44459;
  wire  T_44460;
  wire  T_44461;
  wire  T_44462;
  wire  T_44463;
  wire  T_44464;
  wire  T_44465;
  wire  T_44466;
  wire  T_44467;
  wire  T_44468;
  wire  T_44469;
  wire  T_44470;
  wire  T_44471;
  wire  T_44480;
  wire  T_44481;
  wire  T_44482;
  wire  T_44483;
  wire  T_44484;
  wire  T_44485;
  wire  T_44486;
  wire  T_44487;
  wire  T_44488;
  wire  T_44489;
  wire  T_44490;
  wire  T_44491;
  wire  T_44492;
  wire  T_44493;
  wire  T_44494;
  wire  T_44495;
  wire  T_44496;
  wire  T_44497;
  wire  T_44498;
  wire  T_44499;
  wire  T_44500;
  wire  T_44501;
  wire  T_44502;
  wire  T_44503;
  wire  T_44512;
  wire  T_44513;
  wire  T_44514;
  wire  T_44515;
  wire  T_44516;
  wire  T_44517;
  wire  T_44518;
  wire  T_44519;
  wire  T_44520;
  wire  T_44521;
  wire  T_44522;
  wire  T_44523;
  wire  T_44524;
  wire  T_44525;
  wire  T_44526;
  wire  T_44527;
  wire  T_44528;
  wire  T_44529;
  wire  T_44530;
  wire  T_44531;
  wire  T_44532;
  wire  T_44533;
  wire  T_44534;
  wire  T_44535;
  wire  T_44543;
  wire  T_44544;
  wire  T_44545;
  wire  T_44546;
  wire  T_44547;
  wire  T_44548;
  wire  T_44549;
  wire  T_44550;
  wire  T_44551;
  wire  T_44552;
  wire  T_44553;
  wire  T_44554;
  wire  T_44555;
  wire  T_44556;
  wire  T_44557;
  wire  T_44558;
  wire  T_44559;
  wire  T_44560;
  wire  T_44561;
  wire  T_44562;
  wire  T_44563;
  wire  T_44564;
  wire  T_44565;
  wire  T_44566;
  wire  T_44567;
  wire  T_44575;
  wire  T_44576;
  wire  T_44577;
  wire  T_44578;
  wire  T_44579;
  wire  T_44580;
  wire  T_44581;
  wire  T_44582;
  wire  T_44583;
  wire  T_44584;
  wire  T_44585;
  wire  T_44586;
  wire  T_44587;
  wire  T_44588;
  wire  T_44589;
  wire  T_44590;
  wire  T_44591;
  wire  T_44592;
  wire  T_44593;
  wire  T_44594;
  wire  T_44595;
  wire  T_44596;
  wire  T_44597;
  wire  T_44598;
  wire  T_44599;
  wire  T_44607;
  wire  T_44608;
  wire  T_44609;
  wire  T_44610;
  wire  T_44611;
  wire  T_44612;
  wire  T_44613;
  wire  T_44614;
  wire  T_44615;
  wire  T_44616;
  wire  T_44617;
  wire  T_44618;
  wire  T_44619;
  wire  T_44620;
  wire  T_44621;
  wire  T_44622;
  wire  T_44623;
  wire  T_44624;
  wire  T_44625;
  wire  T_44626;
  wire  T_44627;
  wire  T_44628;
  wire  T_44629;
  wire  T_44630;
  wire  T_44631;
  wire  T_44639;
  wire  T_44640;
  wire  T_44641;
  wire  T_44642;
  wire  T_44643;
  wire  T_44644;
  wire  T_44645;
  wire  T_44646;
  wire  T_44647;
  wire  T_44648;
  wire  T_44649;
  wire  T_44650;
  wire  T_44651;
  wire  T_44652;
  wire  T_44653;
  wire  T_44654;
  wire  T_44655;
  wire  T_44656;
  wire  T_44657;
  wire  T_44658;
  wire  T_44659;
  wire  T_44660;
  wire  T_44661;
  wire  T_44662;
  wire  T_44663;
  wire  T_44670;
  wire  T_44671;
  wire  T_44672;
  wire  T_44673;
  wire  T_44674;
  wire  T_44675;
  wire  T_44676;
  wire  T_44677;
  wire  T_44678;
  wire  T_44679;
  wire  T_44680;
  wire  T_44681;
  wire  T_44682;
  wire  T_44683;
  wire  T_44684;
  wire  T_44685;
  wire  T_44686;
  wire  T_44687;
  wire  T_44688;
  wire  T_44689;
  wire  T_44690;
  wire  T_44691;
  wire  T_44692;
  wire  T_44693;
  wire  T_44694;
  wire  T_44695;
  wire  T_44702;
  wire  T_44703;
  wire  T_44704;
  wire  T_44705;
  wire  T_44706;
  wire  T_44707;
  wire  T_44708;
  wire  T_44709;
  wire  T_44710;
  wire  T_44711;
  wire  T_44712;
  wire  T_44713;
  wire  T_44714;
  wire  T_44715;
  wire  T_44716;
  wire  T_44717;
  wire  T_44718;
  wire  T_44719;
  wire  T_44720;
  wire  T_44721;
  wire  T_44722;
  wire  T_44723;
  wire  T_44724;
  wire  T_44725;
  wire  T_44726;
  wire  T_44727;
  wire  T_44734;
  wire  T_44735;
  wire  T_44736;
  wire  T_44737;
  wire  T_44738;
  wire  T_44739;
  wire  T_44740;
  wire  T_44741;
  wire  T_44742;
  wire  T_44743;
  wire  T_44744;
  wire  T_44745;
  wire  T_44746;
  wire  T_44747;
  wire  T_44748;
  wire  T_44749;
  wire  T_44750;
  wire  T_44751;
  wire  T_44752;
  wire  T_44753;
  wire  T_44754;
  wire  T_44755;
  wire  T_44756;
  wire  T_44757;
  wire  T_44758;
  wire  T_44759;
  wire  T_44766;
  wire  T_44767;
  wire  T_44768;
  wire  T_44769;
  wire  T_44770;
  wire  T_44771;
  wire  T_44772;
  wire  T_44773;
  wire  T_44774;
  wire  T_44775;
  wire  T_44776;
  wire  T_44777;
  wire  T_44778;
  wire  T_44779;
  wire  T_44780;
  wire  T_44781;
  wire  T_44782;
  wire  T_44783;
  wire  T_44784;
  wire  T_44785;
  wire  T_44786;
  wire  T_44787;
  wire  T_44788;
  wire  T_44789;
  wire  T_44790;
  wire  T_44791;
  wire  T_44797;
  wire  T_44798;
  wire  T_44799;
  wire  T_44800;
  wire  T_44801;
  wire  T_44802;
  wire  T_44803;
  wire  T_44804;
  wire  T_44805;
  wire  T_44806;
  wire  T_44807;
  wire  T_44808;
  wire  T_44809;
  wire  T_44810;
  wire  T_44811;
  wire  T_44812;
  wire  T_44813;
  wire  T_44814;
  wire  T_44815;
  wire  T_44816;
  wire  T_44817;
  wire  T_44818;
  wire  T_44819;
  wire  T_44820;
  wire  T_44821;
  wire  T_44822;
  wire  T_44823;
  wire  T_44829;
  wire  T_44830;
  wire  T_44831;
  wire  T_44832;
  wire  T_44833;
  wire  T_44834;
  wire  T_44835;
  wire  T_44836;
  wire  T_44837;
  wire  T_44838;
  wire  T_44839;
  wire  T_44840;
  wire  T_44841;
  wire  T_44842;
  wire  T_44843;
  wire  T_44844;
  wire  T_44845;
  wire  T_44846;
  wire  T_44847;
  wire  T_44848;
  wire  T_44849;
  wire  T_44850;
  wire  T_44851;
  wire  T_44852;
  wire  T_44853;
  wire  T_44854;
  wire  T_44855;
  wire  T_44861;
  wire  T_44862;
  wire  T_44863;
  wire  T_44864;
  wire  T_44865;
  wire  T_44866;
  wire  T_44867;
  wire  T_44868;
  wire  T_44869;
  wire  T_44870;
  wire  T_44871;
  wire  T_44872;
  wire  T_44873;
  wire  T_44874;
  wire  T_44875;
  wire  T_44876;
  wire  T_44877;
  wire  T_44878;
  wire  T_44879;
  wire  T_44880;
  wire  T_44881;
  wire  T_44882;
  wire  T_44883;
  wire  T_44884;
  wire  T_44885;
  wire  T_44886;
  wire  T_44887;
  wire  T_44893;
  wire  T_44894;
  wire  T_44895;
  wire  T_44896;
  wire  T_44897;
  wire  T_44898;
  wire  T_44899;
  wire  T_44900;
  wire  T_44901;
  wire  T_44902;
  wire  T_44903;
  wire  T_44904;
  wire  T_44905;
  wire  T_44906;
  wire  T_44907;
  wire  T_44908;
  wire  T_44909;
  wire  T_44910;
  wire  T_44911;
  wire  T_44912;
  wire  T_44913;
  wire  T_44914;
  wire  T_44915;
  wire  T_44916;
  wire  T_44917;
  wire  T_44918;
  wire  T_44919;
  wire  T_44924;
  wire  T_44925;
  wire  T_44926;
  wire  T_44927;
  wire  T_44928;
  wire  T_44929;
  wire  T_44930;
  wire  T_44931;
  wire  T_44932;
  wire  T_44933;
  wire  T_44934;
  wire  T_44935;
  wire  T_44936;
  wire  T_44937;
  wire  T_44938;
  wire  T_44939;
  wire  T_44940;
  wire  T_44941;
  wire  T_44942;
  wire  T_44943;
  wire  T_44944;
  wire  T_44945;
  wire  T_44946;
  wire  T_44947;
  wire  T_44948;
  wire  T_44949;
  wire  T_44950;
  wire  T_44951;
  wire  T_44956;
  wire  T_44957;
  wire  T_44958;
  wire  T_44959;
  wire  T_44960;
  wire  T_44961;
  wire  T_44962;
  wire  T_44963;
  wire  T_44964;
  wire  T_44965;
  wire  T_44966;
  wire  T_44967;
  wire  T_44968;
  wire  T_44969;
  wire  T_44970;
  wire  T_44971;
  wire  T_44972;
  wire  T_44973;
  wire  T_44974;
  wire  T_44975;
  wire  T_44976;
  wire  T_44977;
  wire  T_44978;
  wire  T_44979;
  wire  T_44980;
  wire  T_44981;
  wire  T_44982;
  wire  T_44983;
  wire  T_44988;
  wire  T_44989;
  wire  T_44990;
  wire  T_44991;
  wire  T_44992;
  wire  T_44993;
  wire  T_44994;
  wire  T_44995;
  wire  T_44996;
  wire  T_44997;
  wire  T_44998;
  wire  T_44999;
  wire  T_45000;
  wire  T_45001;
  wire  T_45002;
  wire  T_45003;
  wire  T_45004;
  wire  T_45005;
  wire  T_45006;
  wire  T_45007;
  wire  T_45008;
  wire  T_45009;
  wire  T_45010;
  wire  T_45011;
  wire  T_45012;
  wire  T_45013;
  wire  T_45014;
  wire  T_45015;
  wire  T_45020;
  wire  T_45021;
  wire  T_45022;
  wire  T_45023;
  wire  T_45024;
  wire  T_45025;
  wire  T_45026;
  wire  T_45027;
  wire  T_45028;
  wire  T_45029;
  wire  T_45030;
  wire  T_45031;
  wire  T_45032;
  wire  T_45033;
  wire  T_45034;
  wire  T_45035;
  wire  T_45036;
  wire  T_45037;
  wire  T_45038;
  wire  T_45039;
  wire  T_45040;
  wire  T_45041;
  wire  T_45042;
  wire  T_45043;
  wire  T_45044;
  wire  T_45045;
  wire  T_45046;
  wire  T_45047;
  wire  T_45051;
  wire  T_45052;
  wire  T_45053;
  wire  T_45054;
  wire  T_45055;
  wire  T_45056;
  wire  T_45057;
  wire  T_45058;
  wire  T_45059;
  wire  T_45060;
  wire  T_45061;
  wire  T_45062;
  wire  T_45063;
  wire  T_45064;
  wire  T_45065;
  wire  T_45066;
  wire  T_45067;
  wire  T_45068;
  wire  T_45069;
  wire  T_45070;
  wire  T_45071;
  wire  T_45072;
  wire  T_45073;
  wire  T_45074;
  wire  T_45075;
  wire  T_45076;
  wire  T_45077;
  wire  T_45078;
  wire  T_45079;
  wire  T_45083;
  wire  T_45084;
  wire  T_45085;
  wire  T_45086;
  wire  T_45087;
  wire  T_45088;
  wire  T_45089;
  wire  T_45090;
  wire  T_45091;
  wire  T_45092;
  wire  T_45093;
  wire  T_45094;
  wire  T_45095;
  wire  T_45096;
  wire  T_45097;
  wire  T_45098;
  wire  T_45099;
  wire  T_45100;
  wire  T_45101;
  wire  T_45102;
  wire  T_45103;
  wire  T_45104;
  wire  T_45105;
  wire  T_45106;
  wire  T_45107;
  wire  T_45108;
  wire  T_45109;
  wire  T_45110;
  wire  T_45111;
  wire  T_45115;
  wire  T_45116;
  wire  T_45117;
  wire  T_45118;
  wire  T_45119;
  wire  T_45120;
  wire  T_45121;
  wire  T_45122;
  wire  T_45123;
  wire  T_45124;
  wire  T_45125;
  wire  T_45126;
  wire  T_45127;
  wire  T_45128;
  wire  T_45129;
  wire  T_45130;
  wire  T_45131;
  wire  T_45132;
  wire  T_45133;
  wire  T_45134;
  wire  T_45135;
  wire  T_45136;
  wire  T_45137;
  wire  T_45138;
  wire  T_45139;
  wire  T_45140;
  wire  T_45141;
  wire  T_45142;
  wire  T_45143;
  wire  T_45147;
  wire  T_45148;
  wire  T_45149;
  wire  T_45150;
  wire  T_45151;
  wire  T_45152;
  wire  T_45153;
  wire  T_45154;
  wire  T_45155;
  wire  T_45156;
  wire  T_45157;
  wire  T_45158;
  wire  T_45159;
  wire  T_45160;
  wire  T_45161;
  wire  T_45162;
  wire  T_45163;
  wire  T_45164;
  wire  T_45165;
  wire  T_45166;
  wire  T_45167;
  wire  T_45168;
  wire  T_45169;
  wire  T_45170;
  wire  T_45171;
  wire  T_45172;
  wire  T_45173;
  wire  T_45174;
  wire  T_45175;
  wire  T_45178;
  wire  T_45179;
  wire  T_45180;
  wire  T_45181;
  wire  T_45182;
  wire  T_45183;
  wire  T_45184;
  wire  T_45185;
  wire  T_45186;
  wire  T_45187;
  wire  T_45188;
  wire  T_45189;
  wire  T_45190;
  wire  T_45191;
  wire  T_45192;
  wire  T_45193;
  wire  T_45194;
  wire  T_45195;
  wire  T_45196;
  wire  T_45197;
  wire  T_45198;
  wire  T_45199;
  wire  T_45200;
  wire  T_45201;
  wire  T_45202;
  wire  T_45203;
  wire  T_45204;
  wire  T_45205;
  wire  T_45206;
  wire  T_45207;
  wire  T_45210;
  wire  T_45211;
  wire  T_45212;
  wire  T_45213;
  wire  T_45214;
  wire  T_45215;
  wire  T_45216;
  wire  T_45217;
  wire  T_45218;
  wire  T_45219;
  wire  T_45220;
  wire  T_45221;
  wire  T_45222;
  wire  T_45223;
  wire  T_45224;
  wire  T_45225;
  wire  T_45226;
  wire  T_45227;
  wire  T_45228;
  wire  T_45229;
  wire  T_45230;
  wire  T_45231;
  wire  T_45232;
  wire  T_45233;
  wire  T_45234;
  wire  T_45235;
  wire  T_45236;
  wire  T_45237;
  wire  T_45238;
  wire  T_45239;
  wire  T_45242;
  wire  T_45243;
  wire  T_45244;
  wire  T_45245;
  wire  T_45246;
  wire  T_45247;
  wire  T_45248;
  wire  T_45249;
  wire  T_45250;
  wire  T_45251;
  wire  T_45252;
  wire  T_45253;
  wire  T_45254;
  wire  T_45255;
  wire  T_45256;
  wire  T_45257;
  wire  T_45258;
  wire  T_45259;
  wire  T_45260;
  wire  T_45261;
  wire  T_45262;
  wire  T_45263;
  wire  T_45264;
  wire  T_45265;
  wire  T_45266;
  wire  T_45267;
  wire  T_45268;
  wire  T_45269;
  wire  T_45270;
  wire  T_45271;
  wire  T_45274;
  wire  T_45275;
  wire  T_45276;
  wire  T_45277;
  wire  T_45278;
  wire  T_45279;
  wire  T_45280;
  wire  T_45281;
  wire  T_45282;
  wire  T_45283;
  wire  T_45284;
  wire  T_45285;
  wire  T_45286;
  wire  T_45287;
  wire  T_45288;
  wire  T_45289;
  wire  T_45290;
  wire  T_45291;
  wire  T_45292;
  wire  T_45293;
  wire  T_45294;
  wire  T_45295;
  wire  T_45296;
  wire  T_45297;
  wire  T_45298;
  wire  T_45299;
  wire  T_45300;
  wire  T_45301;
  wire  T_45302;
  wire  T_45303;
  wire  T_45305;
  wire  T_45306;
  wire  T_45307;
  wire  T_45308;
  wire  T_45309;
  wire  T_45310;
  wire  T_45311;
  wire  T_45312;
  wire  T_45313;
  wire  T_45314;
  wire  T_45315;
  wire  T_45316;
  wire  T_45317;
  wire  T_45318;
  wire  T_45319;
  wire  T_45320;
  wire  T_45321;
  wire  T_45322;
  wire  T_45323;
  wire  T_45324;
  wire  T_45325;
  wire  T_45326;
  wire  T_45327;
  wire  T_45328;
  wire  T_45329;
  wire  T_45330;
  wire  T_45331;
  wire  T_45332;
  wire  T_45333;
  wire  T_45334;
  wire  T_45335;
  wire  T_45337;
  wire  T_45338;
  wire  T_45339;
  wire  T_45340;
  wire  T_45341;
  wire  T_45342;
  wire  T_45343;
  wire  T_45344;
  wire  T_45345;
  wire  T_45346;
  wire  T_45347;
  wire  T_45348;
  wire  T_45349;
  wire  T_45350;
  wire  T_45351;
  wire  T_45352;
  wire  T_45353;
  wire  T_45354;
  wire  T_45355;
  wire  T_45356;
  wire  T_45357;
  wire  T_45358;
  wire  T_45359;
  wire  T_45360;
  wire  T_45361;
  wire  T_45362;
  wire  T_45363;
  wire  T_45364;
  wire  T_45365;
  wire  T_45366;
  wire  T_45367;
  wire  T_45369;
  wire  T_45370;
  wire  T_45371;
  wire  T_45372;
  wire  T_45373;
  wire  T_45374;
  wire  T_45375;
  wire  T_45376;
  wire  T_45377;
  wire  T_45378;
  wire  T_45379;
  wire  T_45380;
  wire  T_45381;
  wire  T_45382;
  wire  T_45383;
  wire  T_45384;
  wire  T_45385;
  wire  T_45386;
  wire  T_45387;
  wire  T_45388;
  wire  T_45389;
  wire  T_45390;
  wire  T_45391;
  wire  T_45392;
  wire  T_45393;
  wire  T_45394;
  wire  T_45395;
  wire  T_45396;
  wire  T_45397;
  wire  T_45398;
  wire  T_45399;
  wire  T_45401;
  wire  T_45402;
  wire  T_45403;
  wire  T_45404;
  wire  T_45405;
  wire  T_45406;
  wire  T_45407;
  wire  T_45408;
  wire  T_45409;
  wire  T_45410;
  wire  T_45411;
  wire  T_45412;
  wire  T_45413;
  wire  T_45414;
  wire  T_45415;
  wire  T_45416;
  wire  T_45417;
  wire  T_45418;
  wire  T_45419;
  wire  T_45420;
  wire  T_45421;
  wire  T_45422;
  wire  T_45423;
  wire  T_45424;
  wire  T_45425;
  wire  T_45426;
  wire  T_45427;
  wire  T_45428;
  wire  T_45429;
  wire  T_45430;
  wire  T_45431;
  wire  T_45473;
  wire  T_45474;
  wire  T_45475;
  wire  T_45476;
  wire  T_45477;
  wire  T_45478;
  wire  T_45479;
  wire  T_45480;
  wire  T_45481;
  wire  T_45482;
  wire  T_45483;
  wire  T_45484;
  wire  T_45485;
  wire  T_45486;
  wire  T_45487;
  wire  T_45488;
  wire  T_45489;
  wire  T_45490;
  wire  T_45491;
  wire  T_45493;
  wire  T_45494;
  wire  T_45495;
  wire  T_45496;
  wire  T_45497;
  wire  T_45498;
  wire  T_45499;
  wire  T_45500;
  wire  T_45501;
  wire  T_45502;
  wire  T_45503;
  wire  T_45504;
  wire  T_45505;
  wire  T_45506;
  wire  T_45507;
  wire  T_45508;
  wire  T_45509;
  wire  T_45510;
  wire  T_45511;
  wire  T_45513;
  wire  T_45514;
  wire  T_45515;
  wire  T_45516;
  wire  T_45517;
  wire  T_45518;
  wire  T_45519;
  wire  T_45520;
  wire  T_45521;
  wire  T_45522;
  wire  T_45523;
  wire  T_45524;
  wire  T_45525;
  wire  T_45526;
  wire  T_45527;
  wire  T_45528;
  wire  T_45529;
  wire  T_45530;
  wire  T_45531;
  wire  T_45533;
  wire  T_45534;
  wire  T_45535;
  wire  T_45536;
  wire  T_45537;
  wire  T_45538;
  wire  T_45539;
  wire  T_45540;
  wire  T_45541;
  wire  T_45542;
  wire  T_45543;
  wire  T_45544;
  wire  T_45545;
  wire  T_45546;
  wire  T_45547;
  wire  T_45548;
  wire  T_45549;
  wire  T_45550;
  wire  T_45551;
  wire  T_45571;
  wire  T_45591;
  wire  T_45611;
  wire  T_45631;
  wire  T_45650;
  wire  T_45651;
  wire  T_45670;
  wire  T_45671;
  wire  T_45690;
  wire  T_45691;
  wire  T_45710;
  wire  T_45711;
  wire  T_45729;
  wire  T_45730;
  wire  T_45731;
  wire  T_45749;
  wire  T_45750;
  wire  T_45751;
  wire  T_45769;
  wire  T_45770;
  wire  T_45771;
  wire  T_45789;
  wire  T_45790;
  wire  T_45791;
  wire  T_45808;
  wire  T_45809;
  wire  T_45810;
  wire  T_45811;
  wire  T_45828;
  wire  T_45829;
  wire  T_45830;
  wire  T_45831;
  wire  T_45848;
  wire  T_45849;
  wire  T_45850;
  wire  T_45851;
  wire  T_45868;
  wire  T_45869;
  wire  T_45870;
  wire  T_45871;
  wire  T_45887;
  wire  T_45888;
  wire  T_45889;
  wire  T_45890;
  wire  T_45891;
  wire  T_45907;
  wire  T_45908;
  wire  T_45909;
  wire  T_45910;
  wire  T_45911;
  wire  T_45927;
  wire  T_45928;
  wire  T_45929;
  wire  T_45930;
  wire  T_45931;
  wire  T_45947;
  wire  T_45948;
  wire  T_45949;
  wire  T_45950;
  wire  T_45951;
  wire  T_45966;
  wire  T_45967;
  wire  T_45968;
  wire  T_45969;
  wire  T_45970;
  wire  T_45971;
  wire  T_45986;
  wire  T_45987;
  wire  T_45988;
  wire  T_45989;
  wire  T_45990;
  wire  T_45991;
  wire  T_46006;
  wire  T_46007;
  wire  T_46008;
  wire  T_46009;
  wire  T_46010;
  wire  T_46011;
  wire  T_46026;
  wire  T_46027;
  wire  T_46028;
  wire  T_46029;
  wire  T_46030;
  wire  T_46031;
  wire  T_46045;
  wire  T_46046;
  wire  T_46047;
  wire  T_46048;
  wire  T_46049;
  wire  T_46050;
  wire  T_46051;
  wire  T_46065;
  wire  T_46066;
  wire  T_46067;
  wire  T_46068;
  wire  T_46069;
  wire  T_46070;
  wire  T_46071;
  wire  T_46085;
  wire  T_46086;
  wire  T_46087;
  wire  T_46088;
  wire  T_46089;
  wire  T_46090;
  wire  T_46091;
  wire  T_46105;
  wire  T_46106;
  wire  T_46107;
  wire  T_46108;
  wire  T_46109;
  wire  T_46110;
  wire  T_46111;
  wire  T_46124;
  wire  T_46125;
  wire  T_46126;
  wire  T_46127;
  wire  T_46128;
  wire  T_46129;
  wire  T_46130;
  wire  T_46131;
  wire  T_46144;
  wire  T_46145;
  wire  T_46146;
  wire  T_46147;
  wire  T_46148;
  wire  T_46149;
  wire  T_46150;
  wire  T_46151;
  wire  T_46164;
  wire  T_46165;
  wire  T_46166;
  wire  T_46167;
  wire  T_46168;
  wire  T_46169;
  wire  T_46170;
  wire  T_46171;
  wire  T_46184;
  wire  T_46185;
  wire  T_46186;
  wire  T_46187;
  wire  T_46188;
  wire  T_46189;
  wire  T_46190;
  wire  T_46191;
  wire  T_46203;
  wire  T_46204;
  wire  T_46205;
  wire  T_46206;
  wire  T_46207;
  wire  T_46208;
  wire  T_46209;
  wire  T_46210;
  wire  T_46211;
  wire  T_46223;
  wire  T_46224;
  wire  T_46225;
  wire  T_46226;
  wire  T_46227;
  wire  T_46228;
  wire  T_46229;
  wire  T_46230;
  wire  T_46231;
  wire  T_46243;
  wire  T_46244;
  wire  T_46245;
  wire  T_46246;
  wire  T_46247;
  wire  T_46248;
  wire  T_46249;
  wire  T_46250;
  wire  T_46251;
  wire  T_46263;
  wire  T_46264;
  wire  T_46265;
  wire  T_46266;
  wire  T_46267;
  wire  T_46268;
  wire  T_46269;
  wire  T_46270;
  wire  T_46271;
  wire  T_46282;
  wire  T_46283;
  wire  T_46284;
  wire  T_46285;
  wire  T_46286;
  wire  T_46287;
  wire  T_46288;
  wire  T_46289;
  wire  T_46290;
  wire  T_46291;
  wire  T_46302;
  wire  T_46303;
  wire  T_46304;
  wire  T_46305;
  wire  T_46306;
  wire  T_46307;
  wire  T_46308;
  wire  T_46309;
  wire  T_46310;
  wire  T_46311;
  wire  T_46322;
  wire  T_46323;
  wire  T_46324;
  wire  T_46325;
  wire  T_46326;
  wire  T_46327;
  wire  T_46328;
  wire  T_46329;
  wire  T_46330;
  wire  T_46331;
  wire  T_46342;
  wire  T_46343;
  wire  T_46344;
  wire  T_46345;
  wire  T_46346;
  wire  T_46347;
  wire  T_46348;
  wire  T_46349;
  wire  T_46350;
  wire  T_46351;
  wire  T_46361;
  wire  T_46362;
  wire  T_46363;
  wire  T_46364;
  wire  T_46365;
  wire  T_46366;
  wire  T_46367;
  wire  T_46368;
  wire  T_46369;
  wire  T_46370;
  wire  T_46371;
  wire  T_46381;
  wire  T_46382;
  wire  T_46383;
  wire  T_46384;
  wire  T_46385;
  wire  T_46386;
  wire  T_46387;
  wire  T_46388;
  wire  T_46389;
  wire  T_46390;
  wire  T_46391;
  wire  T_46401;
  wire  T_46402;
  wire  T_46403;
  wire  T_46404;
  wire  T_46405;
  wire  T_46406;
  wire  T_46407;
  wire  T_46408;
  wire  T_46409;
  wire  T_46410;
  wire  T_46411;
  wire  T_46421;
  wire  T_46422;
  wire  T_46423;
  wire  T_46424;
  wire  T_46425;
  wire  T_46426;
  wire  T_46427;
  wire  T_46428;
  wire  T_46429;
  wire  T_46430;
  wire  T_46431;
  wire  T_46440;
  wire  T_46441;
  wire  T_46442;
  wire  T_46443;
  wire  T_46444;
  wire  T_46445;
  wire  T_46446;
  wire  T_46447;
  wire  T_46448;
  wire  T_46449;
  wire  T_46450;
  wire  T_46451;
  wire  T_46460;
  wire  T_46461;
  wire  T_46462;
  wire  T_46463;
  wire  T_46464;
  wire  T_46465;
  wire  T_46466;
  wire  T_46467;
  wire  T_46468;
  wire  T_46469;
  wire  T_46470;
  wire  T_46471;
  wire  T_46480;
  wire  T_46481;
  wire  T_46482;
  wire  T_46483;
  wire  T_46484;
  wire  T_46485;
  wire  T_46486;
  wire  T_46487;
  wire  T_46488;
  wire  T_46489;
  wire  T_46490;
  wire  T_46491;
  wire  T_46500;
  wire  T_46501;
  wire  T_46502;
  wire  T_46503;
  wire  T_46504;
  wire  T_46505;
  wire  T_46506;
  wire  T_46507;
  wire  T_46508;
  wire  T_46509;
  wire  T_46510;
  wire  T_46511;
  wire  T_46519;
  wire  T_46520;
  wire  T_46521;
  wire  T_46522;
  wire  T_46523;
  wire  T_46524;
  wire  T_46525;
  wire  T_46526;
  wire  T_46527;
  wire  T_46528;
  wire  T_46529;
  wire  T_46530;
  wire  T_46531;
  wire  T_46539;
  wire  T_46540;
  wire  T_46541;
  wire  T_46542;
  wire  T_46543;
  wire  T_46544;
  wire  T_46545;
  wire  T_46546;
  wire  T_46547;
  wire  T_46548;
  wire  T_46549;
  wire  T_46550;
  wire  T_46551;
  wire  T_46559;
  wire  T_46560;
  wire  T_46561;
  wire  T_46562;
  wire  T_46563;
  wire  T_46564;
  wire  T_46565;
  wire  T_46566;
  wire  T_46567;
  wire  T_46568;
  wire  T_46569;
  wire  T_46570;
  wire  T_46571;
  wire  T_46579;
  wire  T_46580;
  wire  T_46581;
  wire  T_46582;
  wire  T_46583;
  wire  T_46584;
  wire  T_46585;
  wire  T_46586;
  wire  T_46587;
  wire  T_46588;
  wire  T_46589;
  wire  T_46590;
  wire  T_46591;
  wire  T_46598;
  wire  T_46599;
  wire  T_46600;
  wire  T_46601;
  wire  T_46602;
  wire  T_46603;
  wire  T_46604;
  wire  T_46605;
  wire  T_46606;
  wire  T_46607;
  wire  T_46608;
  wire  T_46609;
  wire  T_46610;
  wire  T_46611;
  wire  T_46618;
  wire  T_46619;
  wire  T_46620;
  wire  T_46621;
  wire  T_46622;
  wire  T_46623;
  wire  T_46624;
  wire  T_46625;
  wire  T_46626;
  wire  T_46627;
  wire  T_46628;
  wire  T_46629;
  wire  T_46630;
  wire  T_46631;
  wire  T_46638;
  wire  T_46639;
  wire  T_46640;
  wire  T_46641;
  wire  T_46642;
  wire  T_46643;
  wire  T_46644;
  wire  T_46645;
  wire  T_46646;
  wire  T_46647;
  wire  T_46648;
  wire  T_46649;
  wire  T_46650;
  wire  T_46651;
  wire  T_46658;
  wire  T_46659;
  wire  T_46660;
  wire  T_46661;
  wire  T_46662;
  wire  T_46663;
  wire  T_46664;
  wire  T_46665;
  wire  T_46666;
  wire  T_46667;
  wire  T_46668;
  wire  T_46669;
  wire  T_46670;
  wire  T_46671;
  wire  T_46677;
  wire  T_46678;
  wire  T_46679;
  wire  T_46680;
  wire  T_46681;
  wire  T_46682;
  wire  T_46683;
  wire  T_46684;
  wire  T_46685;
  wire  T_46686;
  wire  T_46687;
  wire  T_46688;
  wire  T_46689;
  wire  T_46690;
  wire  T_46691;
  wire  T_46697;
  wire  T_46698;
  wire  T_46699;
  wire  T_46700;
  wire  T_46701;
  wire  T_46702;
  wire  T_46703;
  wire  T_46704;
  wire  T_46705;
  wire  T_46706;
  wire  T_46707;
  wire  T_46708;
  wire  T_46709;
  wire  T_46710;
  wire  T_46711;
  wire  T_46717;
  wire  T_46718;
  wire  T_46719;
  wire  T_46720;
  wire  T_46721;
  wire  T_46722;
  wire  T_46723;
  wire  T_46724;
  wire  T_46725;
  wire  T_46726;
  wire  T_46727;
  wire  T_46728;
  wire  T_46729;
  wire  T_46730;
  wire  T_46731;
  wire  T_46737;
  wire  T_46738;
  wire  T_46739;
  wire  T_46740;
  wire  T_46741;
  wire  T_46742;
  wire  T_46743;
  wire  T_46744;
  wire  T_46745;
  wire  T_46746;
  wire  T_46747;
  wire  T_46748;
  wire  T_46749;
  wire  T_46750;
  wire  T_46751;
  wire  T_46756;
  wire  T_46757;
  wire  T_46758;
  wire  T_46759;
  wire  T_46760;
  wire  T_46761;
  wire  T_46762;
  wire  T_46763;
  wire  T_46764;
  wire  T_46765;
  wire  T_46766;
  wire  T_46767;
  wire  T_46768;
  wire  T_46769;
  wire  T_46770;
  wire  T_46771;
  wire  T_46776;
  wire  T_46777;
  wire  T_46778;
  wire  T_46779;
  wire  T_46780;
  wire  T_46781;
  wire  T_46782;
  wire  T_46783;
  wire  T_46784;
  wire  T_46785;
  wire  T_46786;
  wire  T_46787;
  wire  T_46788;
  wire  T_46789;
  wire  T_46790;
  wire  T_46791;
  wire  T_46796;
  wire  T_46797;
  wire  T_46798;
  wire  T_46799;
  wire  T_46800;
  wire  T_46801;
  wire  T_46802;
  wire  T_46803;
  wire  T_46804;
  wire  T_46805;
  wire  T_46806;
  wire  T_46807;
  wire  T_46808;
  wire  T_46809;
  wire  T_46810;
  wire  T_46811;
  wire  T_46816;
  wire  T_46817;
  wire  T_46818;
  wire  T_46819;
  wire  T_46820;
  wire  T_46821;
  wire  T_46822;
  wire  T_46823;
  wire  T_46824;
  wire  T_46825;
  wire  T_46826;
  wire  T_46827;
  wire  T_46828;
  wire  T_46829;
  wire  T_46830;
  wire  T_46831;
  wire  T_46835;
  wire  T_46836;
  wire  T_46837;
  wire  T_46838;
  wire  T_46839;
  wire  T_46840;
  wire  T_46841;
  wire  T_46842;
  wire  T_46843;
  wire  T_46844;
  wire  T_46845;
  wire  T_46846;
  wire  T_46847;
  wire  T_46848;
  wire  T_46849;
  wire  T_46850;
  wire  T_46851;
  wire  T_46855;
  wire  T_46856;
  wire  T_46857;
  wire  T_46858;
  wire  T_46859;
  wire  T_46860;
  wire  T_46861;
  wire  T_46862;
  wire  T_46863;
  wire  T_46864;
  wire  T_46865;
  wire  T_46866;
  wire  T_46867;
  wire  T_46868;
  wire  T_46869;
  wire  T_46870;
  wire  T_46871;
  wire  T_46875;
  wire  T_46876;
  wire  T_46877;
  wire  T_46878;
  wire  T_46879;
  wire  T_46880;
  wire  T_46881;
  wire  T_46882;
  wire  T_46883;
  wire  T_46884;
  wire  T_46885;
  wire  T_46886;
  wire  T_46887;
  wire  T_46888;
  wire  T_46889;
  wire  T_46890;
  wire  T_46891;
  wire  T_46895;
  wire  T_46896;
  wire  T_46897;
  wire  T_46898;
  wire  T_46899;
  wire  T_46900;
  wire  T_46901;
  wire  T_46902;
  wire  T_46903;
  wire  T_46904;
  wire  T_46905;
  wire  T_46906;
  wire  T_46907;
  wire  T_46908;
  wire  T_46909;
  wire  T_46910;
  wire  T_46911;
  wire  T_46914;
  wire  T_46915;
  wire  T_46916;
  wire  T_46917;
  wire  T_46918;
  wire  T_46919;
  wire  T_46920;
  wire  T_46921;
  wire  T_46922;
  wire  T_46923;
  wire  T_46924;
  wire  T_46925;
  wire  T_46926;
  wire  T_46927;
  wire  T_46928;
  wire  T_46929;
  wire  T_46930;
  wire  T_46931;
  wire  T_46934;
  wire  T_46935;
  wire  T_46936;
  wire  T_46937;
  wire  T_46938;
  wire  T_46939;
  wire  T_46940;
  wire  T_46941;
  wire  T_46942;
  wire  T_46943;
  wire  T_46944;
  wire  T_46945;
  wire  T_46946;
  wire  T_46947;
  wire  T_46948;
  wire  T_46949;
  wire  T_46950;
  wire  T_46951;
  wire  T_46954;
  wire  T_46955;
  wire  T_46956;
  wire  T_46957;
  wire  T_46958;
  wire  T_46959;
  wire  T_46960;
  wire  T_46961;
  wire  T_46962;
  wire  T_46963;
  wire  T_46964;
  wire  T_46965;
  wire  T_46966;
  wire  T_46967;
  wire  T_46968;
  wire  T_46969;
  wire  T_46970;
  wire  T_46971;
  wire  T_46974;
  wire  T_46975;
  wire  T_46976;
  wire  T_46977;
  wire  T_46978;
  wire  T_46979;
  wire  T_46980;
  wire  T_46981;
  wire  T_46982;
  wire  T_46983;
  wire  T_46984;
  wire  T_46985;
  wire  T_46986;
  wire  T_46987;
  wire  T_46988;
  wire  T_46989;
  wire  T_46990;
  wire  T_46991;
  wire  T_46993;
  wire  T_46994;
  wire  T_46995;
  wire  T_46996;
  wire  T_46997;
  wire  T_46998;
  wire  T_46999;
  wire  T_47000;
  wire  T_47001;
  wire  T_47002;
  wire  T_47003;
  wire  T_47004;
  wire  T_47005;
  wire  T_47006;
  wire  T_47007;
  wire  T_47008;
  wire  T_47009;
  wire  T_47010;
  wire  T_47011;
  wire  T_47013;
  wire  T_47014;
  wire  T_47015;
  wire  T_47016;
  wire  T_47017;
  wire  T_47018;
  wire  T_47019;
  wire  T_47020;
  wire  T_47021;
  wire  T_47022;
  wire  T_47023;
  wire  T_47024;
  wire  T_47025;
  wire  T_47026;
  wire  T_47027;
  wire  T_47028;
  wire  T_47029;
  wire  T_47030;
  wire  T_47031;
  wire  T_47033;
  wire  T_47034;
  wire  T_47035;
  wire  T_47036;
  wire  T_47037;
  wire  T_47038;
  wire  T_47039;
  wire  T_47040;
  wire  T_47041;
  wire  T_47042;
  wire  T_47043;
  wire  T_47044;
  wire  T_47045;
  wire  T_47046;
  wire  T_47047;
  wire  T_47048;
  wire  T_47049;
  wire  T_47050;
  wire  T_47051;
  wire  T_47053;
  wire  T_47054;
  wire  T_47055;
  wire  T_47056;
  wire  T_47057;
  wire  T_47058;
  wire  T_47059;
  wire  T_47060;
  wire  T_47061;
  wire  T_47062;
  wire  T_47063;
  wire  T_47064;
  wire  T_47065;
  wire  T_47066;
  wire  T_47067;
  wire  T_47068;
  wire  T_47069;
  wire  T_47070;
  wire  T_47071;
  wire  T_47656_0;
  wire  T_47656_1;
  wire  T_47656_2;
  wire  T_47656_3;
  wire  T_47656_4;
  wire  T_47656_5;
  wire  T_47656_6;
  wire  T_47656_7;
  wire  T_47656_8;
  wire  T_47656_9;
  wire  T_47656_10;
  wire  T_47656_11;
  wire  T_47656_12;
  wire  T_47656_13;
  wire  T_47656_14;
  wire  T_47656_15;
  wire  T_47656_16;
  wire  T_47656_17;
  wire  T_47656_18;
  wire  T_47656_19;
  wire  T_47656_20;
  wire  T_47656_21;
  wire  T_47656_22;
  wire  T_47656_23;
  wire  T_47656_24;
  wire  T_47656_25;
  wire  T_47656_26;
  wire  T_47656_27;
  wire  T_47656_28;
  wire  T_47656_29;
  wire  T_47656_30;
  wire  T_47656_31;
  wire  T_47656_32;
  wire  T_47656_33;
  wire  T_47656_34;
  wire  T_47656_35;
  wire  T_47656_36;
  wire  T_47656_37;
  wire  T_47656_38;
  wire  T_47656_39;
  wire  T_47656_40;
  wire  T_47656_41;
  wire  T_47656_42;
  wire  T_47656_43;
  wire  T_47656_44;
  wire  T_47656_45;
  wire  T_47656_46;
  wire  T_47656_47;
  wire  T_47656_48;
  wire  T_47656_49;
  wire  T_47656_50;
  wire  T_47656_51;
  wire  T_47656_52;
  wire  T_47656_53;
  wire  T_47656_54;
  wire  T_47656_55;
  wire  T_47656_56;
  wire  T_47656_57;
  wire  T_47656_58;
  wire  T_47656_59;
  wire  T_47656_60;
  wire  T_47656_61;
  wire  T_47656_62;
  wire  T_47656_63;
  wire  T_47656_64;
  wire  T_47656_65;
  wire  T_47656_66;
  wire  T_47656_67;
  wire  T_47656_68;
  wire  T_47656_69;
  wire  T_47656_70;
  wire  T_47656_71;
  wire  T_47656_72;
  wire  T_47656_73;
  wire  T_47656_74;
  wire  T_47656_75;
  wire  T_47656_76;
  wire  T_47656_77;
  wire  T_47656_78;
  wire  T_47656_79;
  wire  T_47656_80;
  wire  T_47656_81;
  wire  T_47656_82;
  wire  T_47656_83;
  wire  T_47656_84;
  wire  T_47656_85;
  wire  T_47656_86;
  wire  T_47656_87;
  wire  T_47656_88;
  wire  T_47656_89;
  wire  T_47656_90;
  wire  T_47656_91;
  wire  T_47656_92;
  wire  T_47656_93;
  wire  T_47656_94;
  wire  T_47656_95;
  wire  T_47656_96;
  wire  T_47656_97;
  wire  T_47656_98;
  wire  T_47656_99;
  wire  T_47656_100;
  wire  T_47656_101;
  wire  T_47656_102;
  wire  T_47656_103;
  wire  T_47656_104;
  wire  T_47656_105;
  wire  T_47656_106;
  wire  T_47656_107;
  wire  T_47656_108;
  wire  T_47656_109;
  wire  T_47656_110;
  wire  T_47656_111;
  wire  T_47656_112;
  wire  T_47656_113;
  wire  T_47656_114;
  wire  T_47656_115;
  wire  T_47656_116;
  wire  T_47656_117;
  wire  T_47656_118;
  wire  T_47656_119;
  wire  T_47656_120;
  wire  T_47656_121;
  wire  T_47656_122;
  wire  T_47656_123;
  wire  T_47656_124;
  wire  T_47656_125;
  wire  T_47656_126;
  wire  T_47656_127;
  wire  T_47656_128;
  wire  T_47656_129;
  wire  T_47656_130;
  wire  T_47656_131;
  wire  T_47656_132;
  wire  T_47656_133;
  wire  T_47656_134;
  wire  T_47656_135;
  wire  T_47656_136;
  wire  T_47656_137;
  wire  T_47656_138;
  wire  T_47656_139;
  wire  T_47656_140;
  wire  T_47656_141;
  wire  T_47656_142;
  wire  T_47656_143;
  wire  T_47656_144;
  wire  T_47656_145;
  wire  T_47656_146;
  wire  T_47656_147;
  wire  T_47656_148;
  wire  T_47656_149;
  wire  T_47656_150;
  wire  T_47656_151;
  wire  T_47656_152;
  wire  T_47656_153;
  wire  T_47656_154;
  wire  T_47656_155;
  wire  T_47656_156;
  wire  T_47656_157;
  wire  T_47656_158;
  wire  T_47656_159;
  wire  T_47656_160;
  wire  T_47656_161;
  wire  T_47656_162;
  wire  T_47656_163;
  wire  T_47656_164;
  wire  T_47656_165;
  wire  T_47656_166;
  wire  T_47656_167;
  wire  T_47656_168;
  wire  T_47656_169;
  wire  T_47656_170;
  wire  T_47656_171;
  wire  T_47656_172;
  wire  T_47656_173;
  wire  T_47656_174;
  wire  T_47656_175;
  wire  T_47656_176;
  wire  T_47656_177;
  wire  T_47656_178;
  wire  T_47656_179;
  wire  T_47656_180;
  wire  T_47656_181;
  wire  T_47656_182;
  wire  T_47656_183;
  wire  T_47656_184;
  wire  T_47656_185;
  wire  T_47656_186;
  wire  T_47656_187;
  wire  T_47656_188;
  wire  T_47656_189;
  wire  T_47656_190;
  wire  T_47656_191;
  wire  T_47656_192;
  wire  T_47656_193;
  wire  T_47656_194;
  wire  T_47656_195;
  wire  T_47656_196;
  wire  T_47656_197;
  wire  T_47656_198;
  wire  T_47656_199;
  wire  T_47656_200;
  wire  T_47656_201;
  wire  T_47656_202;
  wire  T_47656_203;
  wire  T_47656_204;
  wire  T_47656_205;
  wire  T_47656_206;
  wire  T_47656_207;
  wire  T_47656_208;
  wire  T_47656_209;
  wire  T_47656_210;
  wire  T_47656_211;
  wire  T_47656_212;
  wire  T_47656_213;
  wire  T_47656_214;
  wire  T_47656_215;
  wire  T_47656_216;
  wire  T_47656_217;
  wire  T_47656_218;
  wire  T_47656_219;
  wire  T_47656_220;
  wire  T_47656_221;
  wire  T_47656_222;
  wire  T_47656_223;
  wire  T_47656_224;
  wire  T_47656_225;
  wire  T_47656_226;
  wire  T_47656_227;
  wire  T_47656_228;
  wire  T_47656_229;
  wire  T_47656_230;
  wire  T_47656_231;
  wire  T_47656_232;
  wire  T_47656_233;
  wire  T_47656_234;
  wire  T_47656_235;
  wire  T_47656_236;
  wire  T_47656_237;
  wire  T_47656_238;
  wire  T_47656_239;
  wire  T_47656_240;
  wire  T_47656_241;
  wire  T_47656_242;
  wire  T_47656_243;
  wire  T_47656_244;
  wire  T_47656_245;
  wire  T_47656_246;
  wire  T_47656_247;
  wire  T_47656_248;
  wire  T_47656_249;
  wire  T_47656_250;
  wire  T_47656_251;
  wire  T_47656_252;
  wire  T_47656_253;
  wire  T_47656_254;
  wire  T_47656_255;
  wire  T_47656_256;
  wire  T_47656_257;
  wire  T_47656_258;
  wire  T_47656_259;
  wire  T_47656_260;
  wire  T_47656_261;
  wire  T_47656_262;
  wire  T_47656_263;
  wire  T_47656_264;
  wire  T_47656_265;
  wire  T_47656_266;
  wire  T_47656_267;
  wire  T_47656_268;
  wire  T_47656_269;
  wire  T_47656_270;
  wire  T_47656_271;
  wire  T_47656_272;
  wire  T_47656_273;
  wire  T_47656_274;
  wire  T_47656_275;
  wire  T_47656_276;
  wire  T_47656_277;
  wire  T_47656_278;
  wire  T_47656_279;
  wire  T_47656_280;
  wire  T_47656_281;
  wire  T_47656_282;
  wire  T_47656_283;
  wire  T_47656_284;
  wire  T_47656_285;
  wire  T_47656_286;
  wire  T_47656_287;
  wire  T_47656_288;
  wire  T_47656_289;
  wire  T_47656_290;
  wire  T_47656_291;
  wire  T_47656_292;
  wire  T_47656_293;
  wire  T_47656_294;
  wire  T_47656_295;
  wire  T_47656_296;
  wire  T_47656_297;
  wire  T_47656_298;
  wire  T_47656_299;
  wire  T_47656_300;
  wire  T_47656_301;
  wire  T_47656_302;
  wire  T_47656_303;
  wire  T_47656_304;
  wire  T_47656_305;
  wire  T_47656_306;
  wire  T_47656_307;
  wire  T_47656_308;
  wire  T_47656_309;
  wire  T_47656_310;
  wire  T_47656_311;
  wire  T_47656_312;
  wire  T_47656_313;
  wire  T_47656_314;
  wire  T_47656_315;
  wire  T_47656_316;
  wire  T_47656_317;
  wire  T_47656_318;
  wire  T_47656_319;
  wire  T_47656_320;
  wire  T_47656_321;
  wire  T_47656_322;
  wire  T_47656_323;
  wire  T_47656_324;
  wire  T_47656_325;
  wire  T_47656_326;
  wire  T_47656_327;
  wire  T_47656_328;
  wire  T_47656_329;
  wire  T_47656_330;
  wire  T_47656_331;
  wire  T_47656_332;
  wire  T_47656_333;
  wire  T_47656_334;
  wire  T_47656_335;
  wire  T_47656_336;
  wire  T_47656_337;
  wire  T_47656_338;
  wire  T_47656_339;
  wire  T_47656_340;
  wire  T_47656_341;
  wire  T_47656_342;
  wire  T_47656_343;
  wire  T_47656_344;
  wire  T_47656_345;
  wire  T_47656_346;
  wire  T_47656_347;
  wire  T_47656_348;
  wire  T_47656_349;
  wire  T_47656_350;
  wire  T_47656_351;
  wire  T_47656_352;
  wire  T_47656_353;
  wire  T_47656_354;
  wire  T_47656_355;
  wire  T_47656_356;
  wire  T_47656_357;
  wire  T_47656_358;
  wire  T_47656_359;
  wire  T_47656_360;
  wire  T_47656_361;
  wire  T_47656_362;
  wire  T_47656_363;
  wire  T_47656_364;
  wire  T_47656_365;
  wire  T_47656_366;
  wire  T_47656_367;
  wire  T_47656_368;
  wire  T_47656_369;
  wire  T_47656_370;
  wire  T_47656_371;
  wire  T_47656_372;
  wire  T_47656_373;
  wire  T_47656_374;
  wire  T_47656_375;
  wire  T_47656_376;
  wire  T_47656_377;
  wire  T_47656_378;
  wire  T_47656_379;
  wire  T_47656_380;
  wire  T_47656_381;
  wire  T_47656_382;
  wire  T_47656_383;
  wire  T_47656_384;
  wire  T_47656_385;
  wire  T_47656_386;
  wire  T_47656_387;
  wire  T_47656_388;
  wire  T_47656_389;
  wire  T_47656_390;
  wire  T_47656_391;
  wire  T_47656_392;
  wire  T_47656_393;
  wire  T_47656_394;
  wire  T_47656_395;
  wire  T_47656_396;
  wire  T_47656_397;
  wire  T_47656_398;
  wire  T_47656_399;
  wire  T_47656_400;
  wire  T_47656_401;
  wire  T_47656_402;
  wire  T_47656_403;
  wire  T_47656_404;
  wire  T_47656_405;
  wire  T_47656_406;
  wire  T_47656_407;
  wire  T_47656_408;
  wire  T_47656_409;
  wire  T_47656_410;
  wire  T_47656_411;
  wire  T_47656_412;
  wire  T_47656_413;
  wire  T_47656_414;
  wire  T_47656_415;
  wire  T_47656_416;
  wire  T_47656_417;
  wire  T_47656_418;
  wire  T_47656_419;
  wire  T_47656_420;
  wire  T_47656_421;
  wire  T_47656_422;
  wire  T_47656_423;
  wire  T_47656_424;
  wire  T_47656_425;
  wire  T_47656_426;
  wire  T_47656_427;
  wire  T_47656_428;
  wire  T_47656_429;
  wire  T_47656_430;
  wire  T_47656_431;
  wire  T_47656_432;
  wire  T_47656_433;
  wire  T_47656_434;
  wire  T_47656_435;
  wire  T_47656_436;
  wire  T_47656_437;
  wire  T_47656_438;
  wire  T_47656_439;
  wire  T_47656_440;
  wire  T_47656_441;
  wire  T_47656_442;
  wire  T_47656_443;
  wire  T_47656_444;
  wire  T_47656_445;
  wire  T_47656_446;
  wire  T_47656_447;
  wire  T_47656_448;
  wire  T_47656_449;
  wire  T_47656_450;
  wire  T_47656_451;
  wire  T_47656_452;
  wire  T_47656_453;
  wire  T_47656_454;
  wire  T_47656_455;
  wire  T_47656_456;
  wire  T_47656_457;
  wire  T_47656_458;
  wire  T_47656_459;
  wire  T_47656_460;
  wire  T_47656_461;
  wire  T_47656_462;
  wire  T_47656_463;
  wire  T_47656_464;
  wire  T_47656_465;
  wire  T_47656_466;
  wire  T_47656_467;
  wire  T_47656_468;
  wire  T_47656_469;
  wire  T_47656_470;
  wire  T_47656_471;
  wire  T_47656_472;
  wire  T_47656_473;
  wire  T_47656_474;
  wire  T_47656_475;
  wire  T_47656_476;
  wire  T_47656_477;
  wire  T_47656_478;
  wire  T_47656_479;
  wire  T_47656_480;
  wire  T_47656_481;
  wire  T_47656_482;
  wire  T_47656_483;
  wire  T_47656_484;
  wire  T_47656_485;
  wire  T_47656_486;
  wire  T_47656_487;
  wire  T_47656_488;
  wire  T_47656_489;
  wire  T_47656_490;
  wire  T_47656_491;
  wire  T_47656_492;
  wire  T_47656_493;
  wire  T_47656_494;
  wire  T_47656_495;
  wire  T_47656_496;
  wire  T_47656_497;
  wire  T_47656_498;
  wire  T_47656_499;
  wire  T_47656_500;
  wire  T_47656_501;
  wire  T_47656_502;
  wire  T_47656_503;
  wire  T_47656_504;
  wire  T_47656_505;
  wire  T_47656_506;
  wire  T_47656_507;
  wire  T_47656_508;
  wire  T_47656_509;
  wire  T_47656_510;
  wire  T_47656_511;
  wire [31:0] T_48687_0;
  wire [31:0] T_48687_1;
  wire [31:0] T_48687_2;
  wire [31:0] T_48687_3;
  wire [31:0] T_48687_4;
  wire [31:0] T_48687_5;
  wire [31:0] T_48687_6;
  wire [31:0] T_48687_7;
  wire [31:0] T_48687_8;
  wire [31:0] T_48687_9;
  wire [31:0] T_48687_10;
  wire [31:0] T_48687_11;
  wire [31:0] T_48687_12;
  wire [31:0] T_48687_13;
  wire [31:0] T_48687_14;
  wire [31:0] T_48687_15;
  wire [31:0] T_48687_16;
  wire [31:0] T_48687_17;
  wire [31:0] T_48687_18;
  wire [31:0] T_48687_19;
  wire [31:0] T_48687_20;
  wire [31:0] T_48687_21;
  wire [31:0] T_48687_22;
  wire [31:0] T_48687_23;
  wire [31:0] T_48687_24;
  wire [31:0] T_48687_25;
  wire [31:0] T_48687_26;
  wire [31:0] T_48687_27;
  wire [31:0] T_48687_28;
  wire [31:0] T_48687_29;
  wire [31:0] T_48687_30;
  wire [31:0] T_48687_31;
  wire [31:0] T_48687_32;
  wire [31:0] T_48687_33;
  wire [31:0] T_48687_34;
  wire [31:0] T_48687_35;
  wire [31:0] T_48687_36;
  wire [31:0] T_48687_37;
  wire [31:0] T_48687_38;
  wire [31:0] T_48687_39;
  wire [31:0] T_48687_40;
  wire [31:0] T_48687_41;
  wire [31:0] T_48687_42;
  wire [31:0] T_48687_43;
  wire [31:0] T_48687_44;
  wire [31:0] T_48687_45;
  wire [31:0] T_48687_46;
  wire [31:0] T_48687_47;
  wire [31:0] T_48687_48;
  wire [31:0] T_48687_49;
  wire [31:0] T_48687_50;
  wire [31:0] T_48687_51;
  wire [31:0] T_48687_52;
  wire [31:0] T_48687_53;
  wire [31:0] T_48687_54;
  wire [31:0] T_48687_55;
  wire [31:0] T_48687_56;
  wire [31:0] T_48687_57;
  wire [31:0] T_48687_58;
  wire [31:0] T_48687_59;
  wire [31:0] T_48687_60;
  wire [31:0] T_48687_61;
  wire [31:0] T_48687_62;
  wire [31:0] T_48687_63;
  wire [31:0] T_48687_64;
  wire [31:0] T_48687_65;
  wire [31:0] T_48687_66;
  wire [31:0] T_48687_67;
  wire [31:0] T_48687_68;
  wire [31:0] T_48687_69;
  wire [31:0] T_48687_70;
  wire [31:0] T_48687_71;
  wire [31:0] T_48687_72;
  wire [31:0] T_48687_73;
  wire [31:0] T_48687_74;
  wire [31:0] T_48687_75;
  wire [31:0] T_48687_76;
  wire [31:0] T_48687_77;
  wire [31:0] T_48687_78;
  wire [31:0] T_48687_79;
  wire [31:0] T_48687_80;
  wire [31:0] T_48687_81;
  wire [31:0] T_48687_82;
  wire [31:0] T_48687_83;
  wire [31:0] T_48687_84;
  wire [31:0] T_48687_85;
  wire [31:0] T_48687_86;
  wire [31:0] T_48687_87;
  wire [31:0] T_48687_88;
  wire [31:0] T_48687_89;
  wire [31:0] T_48687_90;
  wire [31:0] T_48687_91;
  wire [31:0] T_48687_92;
  wire [31:0] T_48687_93;
  wire [31:0] T_48687_94;
  wire [31:0] T_48687_95;
  wire [31:0] T_48687_96;
  wire [31:0] T_48687_97;
  wire [31:0] T_48687_98;
  wire [31:0] T_48687_99;
  wire [31:0] T_48687_100;
  wire [31:0] T_48687_101;
  wire [31:0] T_48687_102;
  wire [31:0] T_48687_103;
  wire [31:0] T_48687_104;
  wire [31:0] T_48687_105;
  wire [31:0] T_48687_106;
  wire [31:0] T_48687_107;
  wire [31:0] T_48687_108;
  wire [31:0] T_48687_109;
  wire [31:0] T_48687_110;
  wire [31:0] T_48687_111;
  wire [31:0] T_48687_112;
  wire [31:0] T_48687_113;
  wire [31:0] T_48687_114;
  wire [31:0] T_48687_115;
  wire [31:0] T_48687_116;
  wire [31:0] T_48687_117;
  wire [31:0] T_48687_118;
  wire [31:0] T_48687_119;
  wire [31:0] T_48687_120;
  wire [31:0] T_48687_121;
  wire [31:0] T_48687_122;
  wire [31:0] T_48687_123;
  wire [31:0] T_48687_124;
  wire [31:0] T_48687_125;
  wire [31:0] T_48687_126;
  wire [31:0] T_48687_127;
  wire [31:0] T_48687_128;
  wire [31:0] T_48687_129;
  wire [31:0] T_48687_130;
  wire [31:0] T_48687_131;
  wire [31:0] T_48687_132;
  wire [31:0] T_48687_133;
  wire [31:0] T_48687_134;
  wire [31:0] T_48687_135;
  wire [31:0] T_48687_136;
  wire [31:0] T_48687_137;
  wire [31:0] T_48687_138;
  wire [31:0] T_48687_139;
  wire [31:0] T_48687_140;
  wire [31:0] T_48687_141;
  wire [31:0] T_48687_142;
  wire [31:0] T_48687_143;
  wire [31:0] T_48687_144;
  wire [31:0] T_48687_145;
  wire [31:0] T_48687_146;
  wire [31:0] T_48687_147;
  wire [31:0] T_48687_148;
  wire [31:0] T_48687_149;
  wire [31:0] T_48687_150;
  wire [31:0] T_48687_151;
  wire [31:0] T_48687_152;
  wire [31:0] T_48687_153;
  wire [31:0] T_48687_154;
  wire [31:0] T_48687_155;
  wire [31:0] T_48687_156;
  wire [31:0] T_48687_157;
  wire [31:0] T_48687_158;
  wire [31:0] T_48687_159;
  wire [31:0] T_48687_160;
  wire [31:0] T_48687_161;
  wire [31:0] T_48687_162;
  wire [31:0] T_48687_163;
  wire [31:0] T_48687_164;
  wire [31:0] T_48687_165;
  wire [31:0] T_48687_166;
  wire [31:0] T_48687_167;
  wire [31:0] T_48687_168;
  wire [31:0] T_48687_169;
  wire [31:0] T_48687_170;
  wire [31:0] T_48687_171;
  wire [31:0] T_48687_172;
  wire [31:0] T_48687_173;
  wire [31:0] T_48687_174;
  wire [31:0] T_48687_175;
  wire [31:0] T_48687_176;
  wire [31:0] T_48687_177;
  wire [31:0] T_48687_178;
  wire [31:0] T_48687_179;
  wire [31:0] T_48687_180;
  wire [31:0] T_48687_181;
  wire [31:0] T_48687_182;
  wire [31:0] T_48687_183;
  wire [31:0] T_48687_184;
  wire [31:0] T_48687_185;
  wire [31:0] T_48687_186;
  wire [31:0] T_48687_187;
  wire [31:0] T_48687_188;
  wire [31:0] T_48687_189;
  wire [31:0] T_48687_190;
  wire [31:0] T_48687_191;
  wire [31:0] T_48687_192;
  wire [31:0] T_48687_193;
  wire [31:0] T_48687_194;
  wire [31:0] T_48687_195;
  wire [31:0] T_48687_196;
  wire [31:0] T_48687_197;
  wire [31:0] T_48687_198;
  wire [31:0] T_48687_199;
  wire [31:0] T_48687_200;
  wire [31:0] T_48687_201;
  wire [31:0] T_48687_202;
  wire [31:0] T_48687_203;
  wire [31:0] T_48687_204;
  wire [31:0] T_48687_205;
  wire [31:0] T_48687_206;
  wire [31:0] T_48687_207;
  wire [31:0] T_48687_208;
  wire [31:0] T_48687_209;
  wire [31:0] T_48687_210;
  wire [31:0] T_48687_211;
  wire [31:0] T_48687_212;
  wire [31:0] T_48687_213;
  wire [31:0] T_48687_214;
  wire [31:0] T_48687_215;
  wire [31:0] T_48687_216;
  wire [31:0] T_48687_217;
  wire [31:0] T_48687_218;
  wire [31:0] T_48687_219;
  wire [31:0] T_48687_220;
  wire [31:0] T_48687_221;
  wire [31:0] T_48687_222;
  wire [31:0] T_48687_223;
  wire [31:0] T_48687_224;
  wire [31:0] T_48687_225;
  wire [31:0] T_48687_226;
  wire [31:0] T_48687_227;
  wire [31:0] T_48687_228;
  wire [31:0] T_48687_229;
  wire [31:0] T_48687_230;
  wire [31:0] T_48687_231;
  wire [31:0] T_48687_232;
  wire [31:0] T_48687_233;
  wire [31:0] T_48687_234;
  wire [31:0] T_48687_235;
  wire [31:0] T_48687_236;
  wire [31:0] T_48687_237;
  wire [31:0] T_48687_238;
  wire [31:0] T_48687_239;
  wire [31:0] T_48687_240;
  wire [31:0] T_48687_241;
  wire [31:0] T_48687_242;
  wire [31:0] T_48687_243;
  wire [31:0] T_48687_244;
  wire [31:0] T_48687_245;
  wire [31:0] T_48687_246;
  wire [31:0] T_48687_247;
  wire [31:0] T_48687_248;
  wire [31:0] T_48687_249;
  wire [31:0] T_48687_250;
  wire [31:0] T_48687_251;
  wire [31:0] T_48687_252;
  wire [31:0] T_48687_253;
  wire [31:0] T_48687_254;
  wire [31:0] T_48687_255;
  wire [31:0] T_48687_256;
  wire [31:0] T_48687_257;
  wire [31:0] T_48687_258;
  wire [31:0] T_48687_259;
  wire [31:0] T_48687_260;
  wire [31:0] T_48687_261;
  wire [31:0] T_48687_262;
  wire [31:0] T_48687_263;
  wire [31:0] T_48687_264;
  wire [31:0] T_48687_265;
  wire [31:0] T_48687_266;
  wire [31:0] T_48687_267;
  wire [31:0] T_48687_268;
  wire [31:0] T_48687_269;
  wire [31:0] T_48687_270;
  wire [31:0] T_48687_271;
  wire [31:0] T_48687_272;
  wire [31:0] T_48687_273;
  wire [31:0] T_48687_274;
  wire [31:0] T_48687_275;
  wire [31:0] T_48687_276;
  wire [31:0] T_48687_277;
  wire [31:0] T_48687_278;
  wire [31:0] T_48687_279;
  wire [31:0] T_48687_280;
  wire [31:0] T_48687_281;
  wire [31:0] T_48687_282;
  wire [31:0] T_48687_283;
  wire [31:0] T_48687_284;
  wire [31:0] T_48687_285;
  wire [31:0] T_48687_286;
  wire [31:0] T_48687_287;
  wire [31:0] T_48687_288;
  wire [31:0] T_48687_289;
  wire [31:0] T_48687_290;
  wire [31:0] T_48687_291;
  wire [31:0] T_48687_292;
  wire [31:0] T_48687_293;
  wire [31:0] T_48687_294;
  wire [31:0] T_48687_295;
  wire [31:0] T_48687_296;
  wire [31:0] T_48687_297;
  wire [31:0] T_48687_298;
  wire [31:0] T_48687_299;
  wire [31:0] T_48687_300;
  wire [31:0] T_48687_301;
  wire [31:0] T_48687_302;
  wire [31:0] T_48687_303;
  wire [31:0] T_48687_304;
  wire [31:0] T_48687_305;
  wire [31:0] T_48687_306;
  wire [31:0] T_48687_307;
  wire [31:0] T_48687_308;
  wire [31:0] T_48687_309;
  wire [31:0] T_48687_310;
  wire [31:0] T_48687_311;
  wire [31:0] T_48687_312;
  wire [31:0] T_48687_313;
  wire [31:0] T_48687_314;
  wire [31:0] T_48687_315;
  wire [31:0] T_48687_316;
  wire [31:0] T_48687_317;
  wire [31:0] T_48687_318;
  wire [31:0] T_48687_319;
  wire [31:0] T_48687_320;
  wire [31:0] T_48687_321;
  wire [31:0] T_48687_322;
  wire [31:0] T_48687_323;
  wire [31:0] T_48687_324;
  wire [31:0] T_48687_325;
  wire [31:0] T_48687_326;
  wire [31:0] T_48687_327;
  wire [31:0] T_48687_328;
  wire [31:0] T_48687_329;
  wire [31:0] T_48687_330;
  wire [31:0] T_48687_331;
  wire [31:0] T_48687_332;
  wire [31:0] T_48687_333;
  wire [31:0] T_48687_334;
  wire [31:0] T_48687_335;
  wire [31:0] T_48687_336;
  wire [31:0] T_48687_337;
  wire [31:0] T_48687_338;
  wire [31:0] T_48687_339;
  wire [31:0] T_48687_340;
  wire [31:0] T_48687_341;
  wire [31:0] T_48687_342;
  wire [31:0] T_48687_343;
  wire [31:0] T_48687_344;
  wire [31:0] T_48687_345;
  wire [31:0] T_48687_346;
  wire [31:0] T_48687_347;
  wire [31:0] T_48687_348;
  wire [31:0] T_48687_349;
  wire [31:0] T_48687_350;
  wire [31:0] T_48687_351;
  wire [31:0] T_48687_352;
  wire [31:0] T_48687_353;
  wire [31:0] T_48687_354;
  wire [31:0] T_48687_355;
  wire [31:0] T_48687_356;
  wire [31:0] T_48687_357;
  wire [31:0] T_48687_358;
  wire [31:0] T_48687_359;
  wire [31:0] T_48687_360;
  wire [31:0] T_48687_361;
  wire [31:0] T_48687_362;
  wire [31:0] T_48687_363;
  wire [31:0] T_48687_364;
  wire [31:0] T_48687_365;
  wire [31:0] T_48687_366;
  wire [31:0] T_48687_367;
  wire [31:0] T_48687_368;
  wire [31:0] T_48687_369;
  wire [31:0] T_48687_370;
  wire [31:0] T_48687_371;
  wire [31:0] T_48687_372;
  wire [31:0] T_48687_373;
  wire [31:0] T_48687_374;
  wire [31:0] T_48687_375;
  wire [31:0] T_48687_376;
  wire [31:0] T_48687_377;
  wire [31:0] T_48687_378;
  wire [31:0] T_48687_379;
  wire [31:0] T_48687_380;
  wire [31:0] T_48687_381;
  wire [31:0] T_48687_382;
  wire [31:0] T_48687_383;
  wire [31:0] T_48687_384;
  wire [31:0] T_48687_385;
  wire [31:0] T_48687_386;
  wire [31:0] T_48687_387;
  wire [31:0] T_48687_388;
  wire [31:0] T_48687_389;
  wire [31:0] T_48687_390;
  wire [31:0] T_48687_391;
  wire [31:0] T_48687_392;
  wire [31:0] T_48687_393;
  wire [31:0] T_48687_394;
  wire [31:0] T_48687_395;
  wire [31:0] T_48687_396;
  wire [31:0] T_48687_397;
  wire [31:0] T_48687_398;
  wire [31:0] T_48687_399;
  wire [31:0] T_48687_400;
  wire [31:0] T_48687_401;
  wire [31:0] T_48687_402;
  wire [31:0] T_48687_403;
  wire [31:0] T_48687_404;
  wire [31:0] T_48687_405;
  wire [31:0] T_48687_406;
  wire [31:0] T_48687_407;
  wire [31:0] T_48687_408;
  wire [31:0] T_48687_409;
  wire [31:0] T_48687_410;
  wire [31:0] T_48687_411;
  wire [31:0] T_48687_412;
  wire [31:0] T_48687_413;
  wire [31:0] T_48687_414;
  wire [31:0] T_48687_415;
  wire [31:0] T_48687_416;
  wire [31:0] T_48687_417;
  wire [31:0] T_48687_418;
  wire [31:0] T_48687_419;
  wire [31:0] T_48687_420;
  wire [31:0] T_48687_421;
  wire [31:0] T_48687_422;
  wire [31:0] T_48687_423;
  wire [31:0] T_48687_424;
  wire [31:0] T_48687_425;
  wire [31:0] T_48687_426;
  wire [31:0] T_48687_427;
  wire [31:0] T_48687_428;
  wire [31:0] T_48687_429;
  wire [31:0] T_48687_430;
  wire [31:0] T_48687_431;
  wire [31:0] T_48687_432;
  wire [31:0] T_48687_433;
  wire [31:0] T_48687_434;
  wire [31:0] T_48687_435;
  wire [31:0] T_48687_436;
  wire [31:0] T_48687_437;
  wire [31:0] T_48687_438;
  wire [31:0] T_48687_439;
  wire [31:0] T_48687_440;
  wire [31:0] T_48687_441;
  wire [31:0] T_48687_442;
  wire [31:0] T_48687_443;
  wire [31:0] T_48687_444;
  wire [31:0] T_48687_445;
  wire [31:0] T_48687_446;
  wire [31:0] T_48687_447;
  wire [31:0] T_48687_448;
  wire [31:0] T_48687_449;
  wire [31:0] T_48687_450;
  wire [31:0] T_48687_451;
  wire [31:0] T_48687_452;
  wire [31:0] T_48687_453;
  wire [31:0] T_48687_454;
  wire [31:0] T_48687_455;
  wire [31:0] T_48687_456;
  wire [31:0] T_48687_457;
  wire [31:0] T_48687_458;
  wire [31:0] T_48687_459;
  wire [31:0] T_48687_460;
  wire [31:0] T_48687_461;
  wire [31:0] T_48687_462;
  wire [31:0] T_48687_463;
  wire [31:0] T_48687_464;
  wire [31:0] T_48687_465;
  wire [31:0] T_48687_466;
  wire [31:0] T_48687_467;
  wire [31:0] T_48687_468;
  wire [31:0] T_48687_469;
  wire [31:0] T_48687_470;
  wire [31:0] T_48687_471;
  wire [31:0] T_48687_472;
  wire [31:0] T_48687_473;
  wire [31:0] T_48687_474;
  wire [31:0] T_48687_475;
  wire [31:0] T_48687_476;
  wire [31:0] T_48687_477;
  wire [31:0] T_48687_478;
  wire [31:0] T_48687_479;
  wire [31:0] T_48687_480;
  wire [31:0] T_48687_481;
  wire [31:0] T_48687_482;
  wire [31:0] T_48687_483;
  wire [31:0] T_48687_484;
  wire [31:0] T_48687_485;
  wire [31:0] T_48687_486;
  wire [31:0] T_48687_487;
  wire [31:0] T_48687_488;
  wire [31:0] T_48687_489;
  wire [31:0] T_48687_490;
  wire [31:0] T_48687_491;
  wire [31:0] T_48687_492;
  wire [31:0] T_48687_493;
  wire [31:0] T_48687_494;
  wire [31:0] T_48687_495;
  wire [31:0] T_48687_496;
  wire [31:0] T_48687_497;
  wire [31:0] T_48687_498;
  wire [31:0] T_48687_499;
  wire [31:0] T_48687_500;
  wire [31:0] T_48687_501;
  wire [31:0] T_48687_502;
  wire [31:0] T_48687_503;
  wire [31:0] T_48687_504;
  wire [31:0] T_48687_505;
  wire [31:0] T_48687_506;
  wire [31:0] T_48687_507;
  wire [31:0] T_48687_508;
  wire [31:0] T_48687_509;
  wire [31:0] T_48687_510;
  wire [31:0] T_48687_511;
  wire  GEN_7;
  wire  GEN_2467;
  wire  GEN_2468;
  wire  GEN_2469;
  wire  GEN_2470;
  wire  GEN_2471;
  wire  GEN_2472;
  wire  GEN_2473;
  wire  GEN_2474;
  wire  GEN_2475;
  wire  GEN_2476;
  wire  GEN_2477;
  wire  GEN_2478;
  wire  GEN_2479;
  wire  GEN_2480;
  wire  GEN_2481;
  wire  GEN_2482;
  wire  GEN_2483;
  wire  GEN_2484;
  wire  GEN_2485;
  wire  GEN_2486;
  wire  GEN_2487;
  wire  GEN_2488;
  wire  GEN_2489;
  wire  GEN_2490;
  wire  GEN_2491;
  wire  GEN_2492;
  wire  GEN_2493;
  wire  GEN_2494;
  wire  GEN_2495;
  wire  GEN_2496;
  wire  GEN_2497;
  wire  GEN_2498;
  wire  GEN_2499;
  wire  GEN_2500;
  wire  GEN_2501;
  wire  GEN_2502;
  wire  GEN_2503;
  wire  GEN_2504;
  wire  GEN_2505;
  wire  GEN_2506;
  wire  GEN_2507;
  wire  GEN_2508;
  wire  GEN_2509;
  wire  GEN_2510;
  wire  GEN_2511;
  wire  GEN_2512;
  wire  GEN_2513;
  wire  GEN_2514;
  wire  GEN_2515;
  wire  GEN_2516;
  wire  GEN_2517;
  wire  GEN_2518;
  wire  GEN_2519;
  wire  GEN_2520;
  wire  GEN_2521;
  wire  GEN_2522;
  wire  GEN_2523;
  wire  GEN_2524;
  wire  GEN_2525;
  wire  GEN_2526;
  wire  GEN_2527;
  wire  GEN_2528;
  wire  GEN_2529;
  wire  GEN_2530;
  wire  GEN_2531;
  wire  GEN_2532;
  wire  GEN_2533;
  wire  GEN_2534;
  wire  GEN_2535;
  wire  GEN_2536;
  wire  GEN_2537;
  wire  GEN_2538;
  wire  GEN_2539;
  wire  GEN_2540;
  wire  GEN_2541;
  wire  GEN_2542;
  wire  GEN_2543;
  wire  GEN_2544;
  wire  GEN_2545;
  wire  GEN_2546;
  wire  GEN_2547;
  wire  GEN_2548;
  wire  GEN_2549;
  wire  GEN_2550;
  wire  GEN_2551;
  wire  GEN_2552;
  wire  GEN_2553;
  wire  GEN_2554;
  wire  GEN_2555;
  wire  GEN_2556;
  wire  GEN_2557;
  wire  GEN_2558;
  wire  GEN_2559;
  wire  GEN_2560;
  wire  GEN_2561;
  wire  GEN_2562;
  wire  GEN_2563;
  wire  GEN_2564;
  wire  GEN_2565;
  wire  GEN_2566;
  wire  GEN_2567;
  wire  GEN_2568;
  wire  GEN_2569;
  wire  GEN_2570;
  wire  GEN_2571;
  wire  GEN_2572;
  wire  GEN_2573;
  wire  GEN_2574;
  wire  GEN_2575;
  wire  GEN_2576;
  wire  GEN_2577;
  wire  GEN_2578;
  wire  GEN_2579;
  wire  GEN_2580;
  wire  GEN_2581;
  wire  GEN_2582;
  wire  GEN_2583;
  wire  GEN_2584;
  wire  GEN_2585;
  wire  GEN_2586;
  wire  GEN_2587;
  wire  GEN_2588;
  wire  GEN_2589;
  wire  GEN_2590;
  wire  GEN_2591;
  wire  GEN_2592;
  wire  GEN_2593;
  wire  GEN_2594;
  wire  GEN_2595;
  wire  GEN_2596;
  wire  GEN_2597;
  wire  GEN_2598;
  wire  GEN_2599;
  wire  GEN_2600;
  wire  GEN_2601;
  wire  GEN_2602;
  wire  GEN_2603;
  wire  GEN_2604;
  wire  GEN_2605;
  wire  GEN_2606;
  wire  GEN_2607;
  wire  GEN_2608;
  wire  GEN_2609;
  wire  GEN_2610;
  wire  GEN_2611;
  wire  GEN_2612;
  wire  GEN_2613;
  wire  GEN_2614;
  wire  GEN_2615;
  wire  GEN_2616;
  wire  GEN_2617;
  wire  GEN_2618;
  wire  GEN_2619;
  wire  GEN_2620;
  wire  GEN_2621;
  wire  GEN_2622;
  wire  GEN_2623;
  wire  GEN_2624;
  wire  GEN_2625;
  wire  GEN_2626;
  wire  GEN_2627;
  wire  GEN_2628;
  wire  GEN_2629;
  wire  GEN_2630;
  wire  GEN_2631;
  wire  GEN_2632;
  wire  GEN_2633;
  wire  GEN_2634;
  wire  GEN_2635;
  wire  GEN_2636;
  wire  GEN_2637;
  wire  GEN_2638;
  wire  GEN_2639;
  wire  GEN_2640;
  wire  GEN_2641;
  wire  GEN_2642;
  wire  GEN_2643;
  wire  GEN_2644;
  wire  GEN_2645;
  wire  GEN_2646;
  wire  GEN_2647;
  wire  GEN_2648;
  wire  GEN_2649;
  wire  GEN_2650;
  wire  GEN_2651;
  wire  GEN_2652;
  wire  GEN_2653;
  wire  GEN_2654;
  wire  GEN_2655;
  wire  GEN_2656;
  wire  GEN_2657;
  wire  GEN_2658;
  wire  GEN_2659;
  wire  GEN_2660;
  wire  GEN_2661;
  wire  GEN_2662;
  wire  GEN_2663;
  wire  GEN_2664;
  wire  GEN_2665;
  wire  GEN_2666;
  wire  GEN_2667;
  wire  GEN_2668;
  wire  GEN_2669;
  wire  GEN_2670;
  wire  GEN_2671;
  wire  GEN_2672;
  wire  GEN_2673;
  wire  GEN_2674;
  wire  GEN_2675;
  wire  GEN_2676;
  wire  GEN_2677;
  wire  GEN_2678;
  wire  GEN_2679;
  wire  GEN_2680;
  wire  GEN_2681;
  wire  GEN_2682;
  wire  GEN_2683;
  wire  GEN_2684;
  wire  GEN_2685;
  wire  GEN_2686;
  wire  GEN_2687;
  wire  GEN_2688;
  wire  GEN_2689;
  wire  GEN_2690;
  wire  GEN_2691;
  wire  GEN_2692;
  wire  GEN_2693;
  wire  GEN_2694;
  wire  GEN_2695;
  wire  GEN_2696;
  wire  GEN_2697;
  wire  GEN_2698;
  wire  GEN_2699;
  wire  GEN_2700;
  wire  GEN_2701;
  wire  GEN_2702;
  wire  GEN_2703;
  wire  GEN_2704;
  wire  GEN_2705;
  wire  GEN_2706;
  wire  GEN_2707;
  wire  GEN_2708;
  wire  GEN_2709;
  wire  GEN_2710;
  wire  GEN_2711;
  wire  GEN_2712;
  wire  GEN_2713;
  wire  GEN_2714;
  wire  GEN_2715;
  wire  GEN_2716;
  wire  GEN_2717;
  wire  GEN_2718;
  wire  GEN_2719;
  wire  GEN_2720;
  wire  GEN_2721;
  wire  GEN_2722;
  wire  GEN_2723;
  wire  GEN_2724;
  wire  GEN_2725;
  wire  GEN_2726;
  wire  GEN_2727;
  wire  GEN_2728;
  wire  GEN_2729;
  wire  GEN_2730;
  wire  GEN_2731;
  wire  GEN_2732;
  wire  GEN_2733;
  wire  GEN_2734;
  wire  GEN_2735;
  wire  GEN_2736;
  wire  GEN_2737;
  wire  GEN_2738;
  wire  GEN_2739;
  wire  GEN_2740;
  wire  GEN_2741;
  wire  GEN_2742;
  wire  GEN_2743;
  wire  GEN_2744;
  wire  GEN_2745;
  wire  GEN_2746;
  wire  GEN_2747;
  wire  GEN_2748;
  wire  GEN_2749;
  wire  GEN_2750;
  wire  GEN_2751;
  wire  GEN_2752;
  wire  GEN_2753;
  wire  GEN_2754;
  wire  GEN_2755;
  wire  GEN_2756;
  wire  GEN_2757;
  wire  GEN_2758;
  wire  GEN_2759;
  wire  GEN_2760;
  wire  GEN_2761;
  wire  GEN_2762;
  wire  GEN_2763;
  wire  GEN_2764;
  wire  GEN_2765;
  wire  GEN_2766;
  wire  GEN_2767;
  wire  GEN_2768;
  wire  GEN_2769;
  wire  GEN_2770;
  wire  GEN_2771;
  wire  GEN_2772;
  wire  GEN_2773;
  wire  GEN_2774;
  wire  GEN_2775;
  wire  GEN_2776;
  wire  GEN_2777;
  wire  GEN_2778;
  wire  GEN_2779;
  wire  GEN_2780;
  wire  GEN_2781;
  wire  GEN_2782;
  wire  GEN_2783;
  wire  GEN_2784;
  wire  GEN_2785;
  wire  GEN_2786;
  wire  GEN_2787;
  wire  GEN_2788;
  wire  GEN_2789;
  wire  GEN_2790;
  wire  GEN_2791;
  wire  GEN_2792;
  wire  GEN_2793;
  wire  GEN_2794;
  wire  GEN_2795;
  wire  GEN_2796;
  wire  GEN_2797;
  wire  GEN_2798;
  wire  GEN_2799;
  wire  GEN_2800;
  wire  GEN_2801;
  wire  GEN_2802;
  wire  GEN_2803;
  wire  GEN_2804;
  wire  GEN_2805;
  wire  GEN_2806;
  wire  GEN_2807;
  wire  GEN_2808;
  wire  GEN_2809;
  wire  GEN_2810;
  wire  GEN_2811;
  wire  GEN_2812;
  wire  GEN_2813;
  wire  GEN_2814;
  wire  GEN_2815;
  wire  GEN_2816;
  wire  GEN_2817;
  wire  GEN_2818;
  wire  GEN_2819;
  wire  GEN_2820;
  wire  GEN_2821;
  wire  GEN_2822;
  wire  GEN_2823;
  wire  GEN_2824;
  wire  GEN_2825;
  wire  GEN_2826;
  wire  GEN_2827;
  wire  GEN_2828;
  wire  GEN_2829;
  wire  GEN_2830;
  wire  GEN_2831;
  wire  GEN_2832;
  wire  GEN_2833;
  wire  GEN_2834;
  wire  GEN_2835;
  wire  GEN_2836;
  wire  GEN_2837;
  wire  GEN_2838;
  wire  GEN_2839;
  wire  GEN_2840;
  wire  GEN_2841;
  wire  GEN_2842;
  wire  GEN_2843;
  wire  GEN_2844;
  wire  GEN_2845;
  wire  GEN_2846;
  wire  GEN_2847;
  wire  GEN_2848;
  wire  GEN_2849;
  wire  GEN_2850;
  wire  GEN_2851;
  wire  GEN_2852;
  wire  GEN_2853;
  wire  GEN_2854;
  wire  GEN_2855;
  wire  GEN_2856;
  wire  GEN_2857;
  wire  GEN_2858;
  wire  GEN_2859;
  wire  GEN_2860;
  wire  GEN_2861;
  wire  GEN_2862;
  wire  GEN_2863;
  wire  GEN_2864;
  wire  GEN_2865;
  wire  GEN_2866;
  wire  GEN_2867;
  wire  GEN_2868;
  wire  GEN_2869;
  wire  GEN_2870;
  wire  GEN_2871;
  wire  GEN_2872;
  wire  GEN_2873;
  wire  GEN_2874;
  wire  GEN_2875;
  wire  GEN_2876;
  wire  GEN_2877;
  wire  GEN_2878;
  wire  GEN_2879;
  wire  GEN_2880;
  wire  GEN_2881;
  wire  GEN_2882;
  wire  GEN_2883;
  wire  GEN_2884;
  wire  GEN_2885;
  wire  GEN_2886;
  wire  GEN_2887;
  wire  GEN_2888;
  wire  GEN_2889;
  wire  GEN_2890;
  wire  GEN_2891;
  wire  GEN_2892;
  wire  GEN_2893;
  wire  GEN_2894;
  wire  GEN_2895;
  wire  GEN_2896;
  wire  GEN_2897;
  wire  GEN_2898;
  wire  GEN_2899;
  wire  GEN_2900;
  wire  GEN_2901;
  wire  GEN_2902;
  wire  GEN_2903;
  wire  GEN_2904;
  wire  GEN_2905;
  wire  GEN_2906;
  wire  GEN_2907;
  wire  GEN_2908;
  wire  GEN_2909;
  wire  GEN_2910;
  wire  GEN_2911;
  wire  GEN_2912;
  wire  GEN_2913;
  wire  GEN_2914;
  wire  GEN_2915;
  wire  GEN_2916;
  wire  GEN_2917;
  wire  GEN_2918;
  wire  GEN_2919;
  wire  GEN_2920;
  wire  GEN_2921;
  wire  GEN_2922;
  wire  GEN_2923;
  wire  GEN_2924;
  wire  GEN_2925;
  wire  GEN_2926;
  wire  GEN_2927;
  wire  GEN_2928;
  wire  GEN_2929;
  wire  GEN_2930;
  wire  GEN_2931;
  wire  GEN_2932;
  wire  GEN_2933;
  wire  GEN_2934;
  wire  GEN_2935;
  wire  GEN_2936;
  wire  GEN_2937;
  wire  GEN_2938;
  wire  GEN_2939;
  wire  GEN_2940;
  wire  GEN_2941;
  wire  GEN_2942;
  wire  GEN_2943;
  wire  GEN_2944;
  wire  GEN_2945;
  wire  GEN_2946;
  wire  GEN_2947;
  wire  GEN_2948;
  wire  GEN_2949;
  wire  GEN_2950;
  wire  GEN_2951;
  wire  GEN_2952;
  wire  GEN_2953;
  wire  GEN_2954;
  wire  GEN_2955;
  wire  GEN_2956;
  wire  GEN_2957;
  wire  GEN_2958;
  wire  GEN_2959;
  wire  GEN_2960;
  wire  GEN_2961;
  wire  GEN_2962;
  wire  GEN_2963;
  wire  GEN_2964;
  wire  GEN_2965;
  wire  GEN_2966;
  wire  GEN_2967;
  wire  GEN_2968;
  wire  GEN_2969;
  wire  GEN_2970;
  wire  GEN_2971;
  wire  GEN_2972;
  wire  GEN_2973;
  wire  GEN_2974;
  wire  GEN_2975;
  wire  GEN_2976;
  wire  GEN_2977;
  wire [31:0] GEN_8;
  wire [31:0] GEN_2978;
  wire [31:0] GEN_2979;
  wire [31:0] GEN_2980;
  wire [31:0] GEN_2981;
  wire [31:0] GEN_2982;
  wire [31:0] GEN_2983;
  wire [31:0] GEN_2984;
  wire [31:0] GEN_2985;
  wire [31:0] GEN_2986;
  wire [31:0] GEN_2987;
  wire [31:0] GEN_2988;
  wire [31:0] GEN_2989;
  wire [31:0] GEN_2990;
  wire [31:0] GEN_2991;
  wire [31:0] GEN_2992;
  wire [31:0] GEN_2993;
  wire [31:0] GEN_2994;
  wire [31:0] GEN_2995;
  wire [31:0] GEN_2996;
  wire [31:0] GEN_2997;
  wire [31:0] GEN_2998;
  wire [31:0] GEN_2999;
  wire [31:0] GEN_3000;
  wire [31:0] GEN_3001;
  wire [31:0] GEN_3002;
  wire [31:0] GEN_3003;
  wire [31:0] GEN_3004;
  wire [31:0] GEN_3005;
  wire [31:0] GEN_3006;
  wire [31:0] GEN_3007;
  wire [31:0] GEN_3008;
  wire [31:0] GEN_3009;
  wire [31:0] GEN_3010;
  wire [31:0] GEN_3011;
  wire [31:0] GEN_3012;
  wire [31:0] GEN_3013;
  wire [31:0] GEN_3014;
  wire [31:0] GEN_3015;
  wire [31:0] GEN_3016;
  wire [31:0] GEN_3017;
  wire [31:0] GEN_3018;
  wire [31:0] GEN_3019;
  wire [31:0] GEN_3020;
  wire [31:0] GEN_3021;
  wire [31:0] GEN_3022;
  wire [31:0] GEN_3023;
  wire [31:0] GEN_3024;
  wire [31:0] GEN_3025;
  wire [31:0] GEN_3026;
  wire [31:0] GEN_3027;
  wire [31:0] GEN_3028;
  wire [31:0] GEN_3029;
  wire [31:0] GEN_3030;
  wire [31:0] GEN_3031;
  wire [31:0] GEN_3032;
  wire [31:0] GEN_3033;
  wire [31:0] GEN_3034;
  wire [31:0] GEN_3035;
  wire [31:0] GEN_3036;
  wire [31:0] GEN_3037;
  wire [31:0] GEN_3038;
  wire [31:0] GEN_3039;
  wire [31:0] GEN_3040;
  wire [31:0] GEN_3041;
  wire [31:0] GEN_3042;
  wire [31:0] GEN_3043;
  wire [31:0] GEN_3044;
  wire [31:0] GEN_3045;
  wire [31:0] GEN_3046;
  wire [31:0] GEN_3047;
  wire [31:0] GEN_3048;
  wire [31:0] GEN_3049;
  wire [31:0] GEN_3050;
  wire [31:0] GEN_3051;
  wire [31:0] GEN_3052;
  wire [31:0] GEN_3053;
  wire [31:0] GEN_3054;
  wire [31:0] GEN_3055;
  wire [31:0] GEN_3056;
  wire [31:0] GEN_3057;
  wire [31:0] GEN_3058;
  wire [31:0] GEN_3059;
  wire [31:0] GEN_3060;
  wire [31:0] GEN_3061;
  wire [31:0] GEN_3062;
  wire [31:0] GEN_3063;
  wire [31:0] GEN_3064;
  wire [31:0] GEN_3065;
  wire [31:0] GEN_3066;
  wire [31:0] GEN_3067;
  wire [31:0] GEN_3068;
  wire [31:0] GEN_3069;
  wire [31:0] GEN_3070;
  wire [31:0] GEN_3071;
  wire [31:0] GEN_3072;
  wire [31:0] GEN_3073;
  wire [31:0] GEN_3074;
  wire [31:0] GEN_3075;
  wire [31:0] GEN_3076;
  wire [31:0] GEN_3077;
  wire [31:0] GEN_3078;
  wire [31:0] GEN_3079;
  wire [31:0] GEN_3080;
  wire [31:0] GEN_3081;
  wire [31:0] GEN_3082;
  wire [31:0] GEN_3083;
  wire [31:0] GEN_3084;
  wire [31:0] GEN_3085;
  wire [31:0] GEN_3086;
  wire [31:0] GEN_3087;
  wire [31:0] GEN_3088;
  wire [31:0] GEN_3089;
  wire [31:0] GEN_3090;
  wire [31:0] GEN_3091;
  wire [31:0] GEN_3092;
  wire [31:0] GEN_3093;
  wire [31:0] GEN_3094;
  wire [31:0] GEN_3095;
  wire [31:0] GEN_3096;
  wire [31:0] GEN_3097;
  wire [31:0] GEN_3098;
  wire [31:0] GEN_3099;
  wire [31:0] GEN_3100;
  wire [31:0] GEN_3101;
  wire [31:0] GEN_3102;
  wire [31:0] GEN_3103;
  wire [31:0] GEN_3104;
  wire [31:0] GEN_3105;
  wire [31:0] GEN_3106;
  wire [31:0] GEN_3107;
  wire [31:0] GEN_3108;
  wire [31:0] GEN_3109;
  wire [31:0] GEN_3110;
  wire [31:0] GEN_3111;
  wire [31:0] GEN_3112;
  wire [31:0] GEN_3113;
  wire [31:0] GEN_3114;
  wire [31:0] GEN_3115;
  wire [31:0] GEN_3116;
  wire [31:0] GEN_3117;
  wire [31:0] GEN_3118;
  wire [31:0] GEN_3119;
  wire [31:0] GEN_3120;
  wire [31:0] GEN_3121;
  wire [31:0] GEN_3122;
  wire [31:0] GEN_3123;
  wire [31:0] GEN_3124;
  wire [31:0] GEN_3125;
  wire [31:0] GEN_3126;
  wire [31:0] GEN_3127;
  wire [31:0] GEN_3128;
  wire [31:0] GEN_3129;
  wire [31:0] GEN_3130;
  wire [31:0] GEN_3131;
  wire [31:0] GEN_3132;
  wire [31:0] GEN_3133;
  wire [31:0] GEN_3134;
  wire [31:0] GEN_3135;
  wire [31:0] GEN_3136;
  wire [31:0] GEN_3137;
  wire [31:0] GEN_3138;
  wire [31:0] GEN_3139;
  wire [31:0] GEN_3140;
  wire [31:0] GEN_3141;
  wire [31:0] GEN_3142;
  wire [31:0] GEN_3143;
  wire [31:0] GEN_3144;
  wire [31:0] GEN_3145;
  wire [31:0] GEN_3146;
  wire [31:0] GEN_3147;
  wire [31:0] GEN_3148;
  wire [31:0] GEN_3149;
  wire [31:0] GEN_3150;
  wire [31:0] GEN_3151;
  wire [31:0] GEN_3152;
  wire [31:0] GEN_3153;
  wire [31:0] GEN_3154;
  wire [31:0] GEN_3155;
  wire [31:0] GEN_3156;
  wire [31:0] GEN_3157;
  wire [31:0] GEN_3158;
  wire [31:0] GEN_3159;
  wire [31:0] GEN_3160;
  wire [31:0] GEN_3161;
  wire [31:0] GEN_3162;
  wire [31:0] GEN_3163;
  wire [31:0] GEN_3164;
  wire [31:0] GEN_3165;
  wire [31:0] GEN_3166;
  wire [31:0] GEN_3167;
  wire [31:0] GEN_3168;
  wire [31:0] GEN_3169;
  wire [31:0] GEN_3170;
  wire [31:0] GEN_3171;
  wire [31:0] GEN_3172;
  wire [31:0] GEN_3173;
  wire [31:0] GEN_3174;
  wire [31:0] GEN_3175;
  wire [31:0] GEN_3176;
  wire [31:0] GEN_3177;
  wire [31:0] GEN_3178;
  wire [31:0] GEN_3179;
  wire [31:0] GEN_3180;
  wire [31:0] GEN_3181;
  wire [31:0] GEN_3182;
  wire [31:0] GEN_3183;
  wire [31:0] GEN_3184;
  wire [31:0] GEN_3185;
  wire [31:0] GEN_3186;
  wire [31:0] GEN_3187;
  wire [31:0] GEN_3188;
  wire [31:0] GEN_3189;
  wire [31:0] GEN_3190;
  wire [31:0] GEN_3191;
  wire [31:0] GEN_3192;
  wire [31:0] GEN_3193;
  wire [31:0] GEN_3194;
  wire [31:0] GEN_3195;
  wire [31:0] GEN_3196;
  wire [31:0] GEN_3197;
  wire [31:0] GEN_3198;
  wire [31:0] GEN_3199;
  wire [31:0] GEN_3200;
  wire [31:0] GEN_3201;
  wire [31:0] GEN_3202;
  wire [31:0] GEN_3203;
  wire [31:0] GEN_3204;
  wire [31:0] GEN_3205;
  wire [31:0] GEN_3206;
  wire [31:0] GEN_3207;
  wire [31:0] GEN_3208;
  wire [31:0] GEN_3209;
  wire [31:0] GEN_3210;
  wire [31:0] GEN_3211;
  wire [31:0] GEN_3212;
  wire [31:0] GEN_3213;
  wire [31:0] GEN_3214;
  wire [31:0] GEN_3215;
  wire [31:0] GEN_3216;
  wire [31:0] GEN_3217;
  wire [31:0] GEN_3218;
  wire [31:0] GEN_3219;
  wire [31:0] GEN_3220;
  wire [31:0] GEN_3221;
  wire [31:0] GEN_3222;
  wire [31:0] GEN_3223;
  wire [31:0] GEN_3224;
  wire [31:0] GEN_3225;
  wire [31:0] GEN_3226;
  wire [31:0] GEN_3227;
  wire [31:0] GEN_3228;
  wire [31:0] GEN_3229;
  wire [31:0] GEN_3230;
  wire [31:0] GEN_3231;
  wire [31:0] GEN_3232;
  wire [31:0] GEN_3233;
  wire [31:0] GEN_3234;
  wire [31:0] GEN_3235;
  wire [31:0] GEN_3236;
  wire [31:0] GEN_3237;
  wire [31:0] GEN_3238;
  wire [31:0] GEN_3239;
  wire [31:0] GEN_3240;
  wire [31:0] GEN_3241;
  wire [31:0] GEN_3242;
  wire [31:0] GEN_3243;
  wire [31:0] GEN_3244;
  wire [31:0] GEN_3245;
  wire [31:0] GEN_3246;
  wire [31:0] GEN_3247;
  wire [31:0] GEN_3248;
  wire [31:0] GEN_3249;
  wire [31:0] GEN_3250;
  wire [31:0] GEN_3251;
  wire [31:0] GEN_3252;
  wire [31:0] GEN_3253;
  wire [31:0] GEN_3254;
  wire [31:0] GEN_3255;
  wire [31:0] GEN_3256;
  wire [31:0] GEN_3257;
  wire [31:0] GEN_3258;
  wire [31:0] GEN_3259;
  wire [31:0] GEN_3260;
  wire [31:0] GEN_3261;
  wire [31:0] GEN_3262;
  wire [31:0] GEN_3263;
  wire [31:0] GEN_3264;
  wire [31:0] GEN_3265;
  wire [31:0] GEN_3266;
  wire [31:0] GEN_3267;
  wire [31:0] GEN_3268;
  wire [31:0] GEN_3269;
  wire [31:0] GEN_3270;
  wire [31:0] GEN_3271;
  wire [31:0] GEN_3272;
  wire [31:0] GEN_3273;
  wire [31:0] GEN_3274;
  wire [31:0] GEN_3275;
  wire [31:0] GEN_3276;
  wire [31:0] GEN_3277;
  wire [31:0] GEN_3278;
  wire [31:0] GEN_3279;
  wire [31:0] GEN_3280;
  wire [31:0] GEN_3281;
  wire [31:0] GEN_3282;
  wire [31:0] GEN_3283;
  wire [31:0] GEN_3284;
  wire [31:0] GEN_3285;
  wire [31:0] GEN_3286;
  wire [31:0] GEN_3287;
  wire [31:0] GEN_3288;
  wire [31:0] GEN_3289;
  wire [31:0] GEN_3290;
  wire [31:0] GEN_3291;
  wire [31:0] GEN_3292;
  wire [31:0] GEN_3293;
  wire [31:0] GEN_3294;
  wire [31:0] GEN_3295;
  wire [31:0] GEN_3296;
  wire [31:0] GEN_3297;
  wire [31:0] GEN_3298;
  wire [31:0] GEN_3299;
  wire [31:0] GEN_3300;
  wire [31:0] GEN_3301;
  wire [31:0] GEN_3302;
  wire [31:0] GEN_3303;
  wire [31:0] GEN_3304;
  wire [31:0] GEN_3305;
  wire [31:0] GEN_3306;
  wire [31:0] GEN_3307;
  wire [31:0] GEN_3308;
  wire [31:0] GEN_3309;
  wire [31:0] GEN_3310;
  wire [31:0] GEN_3311;
  wire [31:0] GEN_3312;
  wire [31:0] GEN_3313;
  wire [31:0] GEN_3314;
  wire [31:0] GEN_3315;
  wire [31:0] GEN_3316;
  wire [31:0] GEN_3317;
  wire [31:0] GEN_3318;
  wire [31:0] GEN_3319;
  wire [31:0] GEN_3320;
  wire [31:0] GEN_3321;
  wire [31:0] GEN_3322;
  wire [31:0] GEN_3323;
  wire [31:0] GEN_3324;
  wire [31:0] GEN_3325;
  wire [31:0] GEN_3326;
  wire [31:0] GEN_3327;
  wire [31:0] GEN_3328;
  wire [31:0] GEN_3329;
  wire [31:0] GEN_3330;
  wire [31:0] GEN_3331;
  wire [31:0] GEN_3332;
  wire [31:0] GEN_3333;
  wire [31:0] GEN_3334;
  wire [31:0] GEN_3335;
  wire [31:0] GEN_3336;
  wire [31:0] GEN_3337;
  wire [31:0] GEN_3338;
  wire [31:0] GEN_3339;
  wire [31:0] GEN_3340;
  wire [31:0] GEN_3341;
  wire [31:0] GEN_3342;
  wire [31:0] GEN_3343;
  wire [31:0] GEN_3344;
  wire [31:0] GEN_3345;
  wire [31:0] GEN_3346;
  wire [31:0] GEN_3347;
  wire [31:0] GEN_3348;
  wire [31:0] GEN_3349;
  wire [31:0] GEN_3350;
  wire [31:0] GEN_3351;
  wire [31:0] GEN_3352;
  wire [31:0] GEN_3353;
  wire [31:0] GEN_3354;
  wire [31:0] GEN_3355;
  wire [31:0] GEN_3356;
  wire [31:0] GEN_3357;
  wire [31:0] GEN_3358;
  wire [31:0] GEN_3359;
  wire [31:0] GEN_3360;
  wire [31:0] GEN_3361;
  wire [31:0] GEN_3362;
  wire [31:0] GEN_3363;
  wire [31:0] GEN_3364;
  wire [31:0] GEN_3365;
  wire [31:0] GEN_3366;
  wire [31:0] GEN_3367;
  wire [31:0] GEN_3368;
  wire [31:0] GEN_3369;
  wire [31:0] GEN_3370;
  wire [31:0] GEN_3371;
  wire [31:0] GEN_3372;
  wire [31:0] GEN_3373;
  wire [31:0] GEN_3374;
  wire [31:0] GEN_3375;
  wire [31:0] GEN_3376;
  wire [31:0] GEN_3377;
  wire [31:0] GEN_3378;
  wire [31:0] GEN_3379;
  wire [31:0] GEN_3380;
  wire [31:0] GEN_3381;
  wire [31:0] GEN_3382;
  wire [31:0] GEN_3383;
  wire [31:0] GEN_3384;
  wire [31:0] GEN_3385;
  wire [31:0] GEN_3386;
  wire [31:0] GEN_3387;
  wire [31:0] GEN_3388;
  wire [31:0] GEN_3389;
  wire [31:0] GEN_3390;
  wire [31:0] GEN_3391;
  wire [31:0] GEN_3392;
  wire [31:0] GEN_3393;
  wire [31:0] GEN_3394;
  wire [31:0] GEN_3395;
  wire [31:0] GEN_3396;
  wire [31:0] GEN_3397;
  wire [31:0] GEN_3398;
  wire [31:0] GEN_3399;
  wire [31:0] GEN_3400;
  wire [31:0] GEN_3401;
  wire [31:0] GEN_3402;
  wire [31:0] GEN_3403;
  wire [31:0] GEN_3404;
  wire [31:0] GEN_3405;
  wire [31:0] GEN_3406;
  wire [31:0] GEN_3407;
  wire [31:0] GEN_3408;
  wire [31:0] GEN_3409;
  wire [31:0] GEN_3410;
  wire [31:0] GEN_3411;
  wire [31:0] GEN_3412;
  wire [31:0] GEN_3413;
  wire [31:0] GEN_3414;
  wire [31:0] GEN_3415;
  wire [31:0] GEN_3416;
  wire [31:0] GEN_3417;
  wire [31:0] GEN_3418;
  wire [31:0] GEN_3419;
  wire [31:0] GEN_3420;
  wire [31:0] GEN_3421;
  wire [31:0] GEN_3422;
  wire [31:0] GEN_3423;
  wire [31:0] GEN_3424;
  wire [31:0] GEN_3425;
  wire [31:0] GEN_3426;
  wire [31:0] GEN_3427;
  wire [31:0] GEN_3428;
  wire [31:0] GEN_3429;
  wire [31:0] GEN_3430;
  wire [31:0] GEN_3431;
  wire [31:0] GEN_3432;
  wire [31:0] GEN_3433;
  wire [31:0] GEN_3434;
  wire [31:0] GEN_3435;
  wire [31:0] GEN_3436;
  wire [31:0] GEN_3437;
  wire [31:0] GEN_3438;
  wire [31:0] GEN_3439;
  wire [31:0] GEN_3440;
  wire [31:0] GEN_3441;
  wire [31:0] GEN_3442;
  wire [31:0] GEN_3443;
  wire [31:0] GEN_3444;
  wire [31:0] GEN_3445;
  wire [31:0] GEN_3446;
  wire [31:0] GEN_3447;
  wire [31:0] GEN_3448;
  wire [31:0] GEN_3449;
  wire [31:0] GEN_3450;
  wire [31:0] GEN_3451;
  wire [31:0] GEN_3452;
  wire [31:0] GEN_3453;
  wire [31:0] GEN_3454;
  wire [31:0] GEN_3455;
  wire [31:0] GEN_3456;
  wire [31:0] GEN_3457;
  wire [31:0] GEN_3458;
  wire [31:0] GEN_3459;
  wire [31:0] GEN_3460;
  wire [31:0] GEN_3461;
  wire [31:0] GEN_3462;
  wire [31:0] GEN_3463;
  wire [31:0] GEN_3464;
  wire [31:0] GEN_3465;
  wire [31:0] GEN_3466;
  wire [31:0] GEN_3467;
  wire [31:0] GEN_3468;
  wire [31:0] GEN_3469;
  wire [31:0] GEN_3470;
  wire [31:0] GEN_3471;
  wire [31:0] GEN_3472;
  wire [31:0] GEN_3473;
  wire [31:0] GEN_3474;
  wire [31:0] GEN_3475;
  wire [31:0] GEN_3476;
  wire [31:0] GEN_3477;
  wire [31:0] GEN_3478;
  wire [31:0] GEN_3479;
  wire [31:0] GEN_3480;
  wire [31:0] GEN_3481;
  wire [31:0] GEN_3482;
  wire [31:0] GEN_3483;
  wire [31:0] GEN_3484;
  wire [31:0] GEN_3485;
  wire [31:0] GEN_3486;
  wire [31:0] GEN_3487;
  wire [31:0] GEN_3488;
  wire [31:0] T_49204;
  wire [1:0] T_49205;
  wire [4:0] T_49207;
  wire [2:0] T_49208;
  wire [2:0] T_49219_opcode;
  wire [1:0] T_49219_param;
  wire [2:0] T_49219_size;
  wire [4:0] T_49219_source;
  wire  T_49219_sink;
  wire [1:0] T_49219_addr_lo;
  wire [31:0] T_49219_data;
  wire  T_49219_error;
  wire [2:0] GEN_60 = 3'b0;
  reg [31:0] GEN_3876;
  wire [1:0] GEN_91 = 2'b0;
  reg [31:0] GEN_3877;
  wire [2:0] GEN_143 = 3'b0;
  reg [31:0] GEN_3878;
  wire [4:0] GEN_364 = 5'b0;
  reg [31:0] GEN_3879;
  wire [27:0] GEN_3714 = 28'b0;
  reg [31:0] GEN_3880;
  wire [3:0] GEN_3715 = 4'b0;
  reg [31:0] GEN_3881;
  wire [31:0] GEN_3716 = 32'b0;
  reg [31:0] GEN_3882;
  sirv_LevelGateway u_LevelGateway_51 (
    .clock(LevelGateway_51_clock),
    .reset(LevelGateway_51_reset),
    .io_interrupt(LevelGateway_51_io_interrupt),
    .io_plic_valid(LevelGateway_51_io_plic_valid),
    .io_plic_ready(LevelGateway_51_io_plic_ready),
    .io_plic_complete(LevelGateway_51_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_1_1 (
    .clock(LevelGateway_1_1_clock),
    .reset(LevelGateway_1_1_reset),
    .io_interrupt(LevelGateway_1_1_io_interrupt),
    .io_plic_valid(LevelGateway_1_1_io_plic_valid),
    .io_plic_ready(LevelGateway_1_1_io_plic_ready),
    .io_plic_complete(LevelGateway_1_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_2_1 (
    .clock(LevelGateway_2_1_clock),
    .reset(LevelGateway_2_1_reset),
    .io_interrupt(LevelGateway_2_1_io_interrupt),
    .io_plic_valid(LevelGateway_2_1_io_plic_valid),
    .io_plic_ready(LevelGateway_2_1_io_plic_ready),
    .io_plic_complete(LevelGateway_2_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_3_1 (
    .clock(LevelGateway_3_1_clock),
    .reset(LevelGateway_3_1_reset),
    .io_interrupt(LevelGateway_3_1_io_interrupt),
    .io_plic_valid(LevelGateway_3_1_io_plic_valid),
    .io_plic_ready(LevelGateway_3_1_io_plic_ready),
    .io_plic_complete(LevelGateway_3_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_4_1 (
    .clock(LevelGateway_4_1_clock),
    .reset(LevelGateway_4_1_reset),
    .io_interrupt(LevelGateway_4_1_io_interrupt),
    .io_plic_valid(LevelGateway_4_1_io_plic_valid),
    .io_plic_ready(LevelGateway_4_1_io_plic_ready),
    .io_plic_complete(LevelGateway_4_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_5_1 (
    .clock(LevelGateway_5_1_clock),
    .reset(LevelGateway_5_1_reset),
    .io_interrupt(LevelGateway_5_1_io_interrupt),
    .io_plic_valid(LevelGateway_5_1_io_plic_valid),
    .io_plic_ready(LevelGateway_5_1_io_plic_ready),
    .io_plic_complete(LevelGateway_5_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_6_1 (
    .clock(LevelGateway_6_1_clock),
    .reset(LevelGateway_6_1_reset),
    .io_interrupt(LevelGateway_6_1_io_interrupt),
    .io_plic_valid(LevelGateway_6_1_io_plic_valid),
    .io_plic_ready(LevelGateway_6_1_io_plic_ready),
    .io_plic_complete(LevelGateway_6_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_7_1 (
    .clock(LevelGateway_7_1_clock),
    .reset(LevelGateway_7_1_reset),
    .io_interrupt(LevelGateway_7_1_io_interrupt),
    .io_plic_valid(LevelGateway_7_1_io_plic_valid),
    .io_plic_ready(LevelGateway_7_1_io_plic_ready),
    .io_plic_complete(LevelGateway_7_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_8_1 (
    .clock(LevelGateway_8_1_clock),
    .reset(LevelGateway_8_1_reset),
    .io_interrupt(LevelGateway_8_1_io_interrupt),
    .io_plic_valid(LevelGateway_8_1_io_plic_valid),
    .io_plic_ready(LevelGateway_8_1_io_plic_ready),
    .io_plic_complete(LevelGateway_8_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_9_1 (
    .clock(LevelGateway_9_1_clock),
    .reset(LevelGateway_9_1_reset),
    .io_interrupt(LevelGateway_9_1_io_interrupt),
    .io_plic_valid(LevelGateway_9_1_io_plic_valid),
    .io_plic_ready(LevelGateway_9_1_io_plic_ready),
    .io_plic_complete(LevelGateway_9_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_10_1 (
    .clock(LevelGateway_10_1_clock),
    .reset(LevelGateway_10_1_reset),
    .io_interrupt(LevelGateway_10_1_io_interrupt),
    .io_plic_valid(LevelGateway_10_1_io_plic_valid),
    .io_plic_ready(LevelGateway_10_1_io_plic_ready),
    .io_plic_complete(LevelGateway_10_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_11_1 (
    .clock(LevelGateway_11_1_clock),
    .reset(LevelGateway_11_1_reset),
    .io_interrupt(LevelGateway_11_1_io_interrupt),
    .io_plic_valid(LevelGateway_11_1_io_plic_valid),
    .io_plic_ready(LevelGateway_11_1_io_plic_ready),
    .io_plic_complete(LevelGateway_11_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_12_1 (
    .clock(LevelGateway_12_1_clock),
    .reset(LevelGateway_12_1_reset),
    .io_interrupt(LevelGateway_12_1_io_interrupt),
    .io_plic_valid(LevelGateway_12_1_io_plic_valid),
    .io_plic_ready(LevelGateway_12_1_io_plic_ready),
    .io_plic_complete(LevelGateway_12_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_13_1 (
    .clock(LevelGateway_13_1_clock),
    .reset(LevelGateway_13_1_reset),
    .io_interrupt(LevelGateway_13_1_io_interrupt),
    .io_plic_valid(LevelGateway_13_1_io_plic_valid),
    .io_plic_ready(LevelGateway_13_1_io_plic_ready),
    .io_plic_complete(LevelGateway_13_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_14_1 (
    .clock(LevelGateway_14_1_clock),
    .reset(LevelGateway_14_1_reset),
    .io_interrupt(LevelGateway_14_1_io_interrupt),
    .io_plic_valid(LevelGateway_14_1_io_plic_valid),
    .io_plic_ready(LevelGateway_14_1_io_plic_ready),
    .io_plic_complete(LevelGateway_14_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_15_1 (
    .clock(LevelGateway_15_1_clock),
    .reset(LevelGateway_15_1_reset),
    .io_interrupt(LevelGateway_15_1_io_interrupt),
    .io_plic_valid(LevelGateway_15_1_io_plic_valid),
    .io_plic_ready(LevelGateway_15_1_io_plic_ready),
    .io_plic_complete(LevelGateway_15_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_16_1 (
    .clock(LevelGateway_16_1_clock),
    .reset(LevelGateway_16_1_reset),
    .io_interrupt(LevelGateway_16_1_io_interrupt),
    .io_plic_valid(LevelGateway_16_1_io_plic_valid),
    .io_plic_ready(LevelGateway_16_1_io_plic_ready),
    .io_plic_complete(LevelGateway_16_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_17_1 (
    .clock(LevelGateway_17_1_clock),
    .reset(LevelGateway_17_1_reset),
    .io_interrupt(LevelGateway_17_1_io_interrupt),
    .io_plic_valid(LevelGateway_17_1_io_plic_valid),
    .io_plic_ready(LevelGateway_17_1_io_plic_ready),
    .io_plic_complete(LevelGateway_17_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_18_1 (
    .clock(LevelGateway_18_1_clock),
    .reset(LevelGateway_18_1_reset),
    .io_interrupt(LevelGateway_18_1_io_interrupt),
    .io_plic_valid(LevelGateway_18_1_io_plic_valid),
    .io_plic_ready(LevelGateway_18_1_io_plic_ready),
    .io_plic_complete(LevelGateway_18_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_19_1 (
    .clock(LevelGateway_19_1_clock),
    .reset(LevelGateway_19_1_reset),
    .io_interrupt(LevelGateway_19_1_io_interrupt),
    .io_plic_valid(LevelGateway_19_1_io_plic_valid),
    .io_plic_ready(LevelGateway_19_1_io_plic_ready),
    .io_plic_complete(LevelGateway_19_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_20_1 (
    .clock(LevelGateway_20_1_clock),
    .reset(LevelGateway_20_1_reset),
    .io_interrupt(LevelGateway_20_1_io_interrupt),
    .io_plic_valid(LevelGateway_20_1_io_plic_valid),
    .io_plic_ready(LevelGateway_20_1_io_plic_ready),
    .io_plic_complete(LevelGateway_20_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_21_1 (
    .clock(LevelGateway_21_1_clock),
    .reset(LevelGateway_21_1_reset),
    .io_interrupt(LevelGateway_21_1_io_interrupt),
    .io_plic_valid(LevelGateway_21_1_io_plic_valid),
    .io_plic_ready(LevelGateway_21_1_io_plic_ready),
    .io_plic_complete(LevelGateway_21_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_22_1 (
    .clock(LevelGateway_22_1_clock),
    .reset(LevelGateway_22_1_reset),
    .io_interrupt(LevelGateway_22_1_io_interrupt),
    .io_plic_valid(LevelGateway_22_1_io_plic_valid),
    .io_plic_ready(LevelGateway_22_1_io_plic_ready),
    .io_plic_complete(LevelGateway_22_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_23_1 (
    .clock(LevelGateway_23_1_clock),
    .reset(LevelGateway_23_1_reset),
    .io_interrupt(LevelGateway_23_1_io_interrupt),
    .io_plic_valid(LevelGateway_23_1_io_plic_valid),
    .io_plic_ready(LevelGateway_23_1_io_plic_ready),
    .io_plic_complete(LevelGateway_23_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_24_1 (
    .clock(LevelGateway_24_1_clock),
    .reset(LevelGateway_24_1_reset),
    .io_interrupt(LevelGateway_24_1_io_interrupt),
    .io_plic_valid(LevelGateway_24_1_io_plic_valid),
    .io_plic_ready(LevelGateway_24_1_io_plic_ready),
    .io_plic_complete(LevelGateway_24_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_25_1 (
    .clock(LevelGateway_25_1_clock),
    .reset(LevelGateway_25_1_reset),
    .io_interrupt(LevelGateway_25_1_io_interrupt),
    .io_plic_valid(LevelGateway_25_1_io_plic_valid),
    .io_plic_ready(LevelGateway_25_1_io_plic_ready),
    .io_plic_complete(LevelGateway_25_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_26_1 (
    .clock(LevelGateway_26_1_clock),
    .reset(LevelGateway_26_1_reset),
    .io_interrupt(LevelGateway_26_1_io_interrupt),
    .io_plic_valid(LevelGateway_26_1_io_plic_valid),
    .io_plic_ready(LevelGateway_26_1_io_plic_ready),
    .io_plic_complete(LevelGateway_26_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_27_1 (
    .clock(LevelGateway_27_1_clock),
    .reset(LevelGateway_27_1_reset),
    .io_interrupt(LevelGateway_27_1_io_interrupt),
    .io_plic_valid(LevelGateway_27_1_io_plic_valid),
    .io_plic_ready(LevelGateway_27_1_io_plic_ready),
    .io_plic_complete(LevelGateway_27_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_28_1 (
    .clock(LevelGateway_28_1_clock),
    .reset(LevelGateway_28_1_reset),
    .io_interrupt(LevelGateway_28_1_io_interrupt),
    .io_plic_valid(LevelGateway_28_1_io_plic_valid),
    .io_plic_ready(LevelGateway_28_1_io_plic_ready),
    .io_plic_complete(LevelGateway_28_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_29_1 (
    .clock(LevelGateway_29_1_clock),
    .reset(LevelGateway_29_1_reset),
    .io_interrupt(LevelGateway_29_1_io_interrupt),
    .io_plic_valid(LevelGateway_29_1_io_plic_valid),
    .io_plic_ready(LevelGateway_29_1_io_plic_ready),
    .io_plic_complete(LevelGateway_29_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_30_1 (
    .clock(LevelGateway_30_1_clock),
    .reset(LevelGateway_30_1_reset),
    .io_interrupt(LevelGateway_30_1_io_interrupt),
    .io_plic_valid(LevelGateway_30_1_io_plic_valid),
    .io_plic_ready(LevelGateway_30_1_io_plic_ready),
    .io_plic_complete(LevelGateway_30_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_31_1 (
    .clock(LevelGateway_31_1_clock),
    .reset(LevelGateway_31_1_reset),
    .io_interrupt(LevelGateway_31_1_io_interrupt),
    .io_plic_valid(LevelGateway_31_1_io_plic_valid),
    .io_plic_ready(LevelGateway_31_1_io_plic_ready),
    .io_plic_complete(LevelGateway_31_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_32_1 (
    .clock(LevelGateway_32_1_clock),
    .reset(LevelGateway_32_1_reset),
    .io_interrupt(LevelGateway_32_1_io_interrupt),
    .io_plic_valid(LevelGateway_32_1_io_plic_valid),
    .io_plic_ready(LevelGateway_32_1_io_plic_ready),
    .io_plic_complete(LevelGateway_32_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_33_1 (
    .clock(LevelGateway_33_1_clock),
    .reset(LevelGateway_33_1_reset),
    .io_interrupt(LevelGateway_33_1_io_interrupt),
    .io_plic_valid(LevelGateway_33_1_io_plic_valid),
    .io_plic_ready(LevelGateway_33_1_io_plic_ready),
    .io_plic_complete(LevelGateway_33_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_34_1 (
    .clock(LevelGateway_34_1_clock),
    .reset(LevelGateway_34_1_reset),
    .io_interrupt(LevelGateway_34_1_io_interrupt),
    .io_plic_valid(LevelGateway_34_1_io_plic_valid),
    .io_plic_ready(LevelGateway_34_1_io_plic_ready),
    .io_plic_complete(LevelGateway_34_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_35_1 (
    .clock(LevelGateway_35_1_clock),
    .reset(LevelGateway_35_1_reset),
    .io_interrupt(LevelGateway_35_1_io_interrupt),
    .io_plic_valid(LevelGateway_35_1_io_plic_valid),
    .io_plic_ready(LevelGateway_35_1_io_plic_ready),
    .io_plic_complete(LevelGateway_35_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_36_1 (
    .clock(LevelGateway_36_1_clock),
    .reset(LevelGateway_36_1_reset),
    .io_interrupt(LevelGateway_36_1_io_interrupt),
    .io_plic_valid(LevelGateway_36_1_io_plic_valid),
    .io_plic_ready(LevelGateway_36_1_io_plic_ready),
    .io_plic_complete(LevelGateway_36_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_37_1 (
    .clock(LevelGateway_37_1_clock),
    .reset(LevelGateway_37_1_reset),
    .io_interrupt(LevelGateway_37_1_io_interrupt),
    .io_plic_valid(LevelGateway_37_1_io_plic_valid),
    .io_plic_ready(LevelGateway_37_1_io_plic_ready),
    .io_plic_complete(LevelGateway_37_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_38_1 (
    .clock(LevelGateway_38_1_clock),
    .reset(LevelGateway_38_1_reset),
    .io_interrupt(LevelGateway_38_1_io_interrupt),
    .io_plic_valid(LevelGateway_38_1_io_plic_valid),
    .io_plic_ready(LevelGateway_38_1_io_plic_ready),
    .io_plic_complete(LevelGateway_38_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_39_1 (
    .clock(LevelGateway_39_1_clock),
    .reset(LevelGateway_39_1_reset),
    .io_interrupt(LevelGateway_39_1_io_interrupt),
    .io_plic_valid(LevelGateway_39_1_io_plic_valid),
    .io_plic_ready(LevelGateway_39_1_io_plic_ready),
    .io_plic_complete(LevelGateway_39_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_40_1 (
    .clock(LevelGateway_40_1_clock),
    .reset(LevelGateway_40_1_reset),
    .io_interrupt(LevelGateway_40_1_io_interrupt),
    .io_plic_valid(LevelGateway_40_1_io_plic_valid),
    .io_plic_ready(LevelGateway_40_1_io_plic_ready),
    .io_plic_complete(LevelGateway_40_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_41_1 (
    .clock(LevelGateway_41_1_clock),
    .reset(LevelGateway_41_1_reset),
    .io_interrupt(LevelGateway_41_1_io_interrupt),
    .io_plic_valid(LevelGateway_41_1_io_plic_valid),
    .io_plic_ready(LevelGateway_41_1_io_plic_ready),
    .io_plic_complete(LevelGateway_41_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_42_1 (
    .clock(LevelGateway_42_1_clock),
    .reset(LevelGateway_42_1_reset),
    .io_interrupt(LevelGateway_42_1_io_interrupt),
    .io_plic_valid(LevelGateway_42_1_io_plic_valid),
    .io_plic_ready(LevelGateway_42_1_io_plic_ready),
    .io_plic_complete(LevelGateway_42_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_43_1 (
    .clock(LevelGateway_43_1_clock),
    .reset(LevelGateway_43_1_reset),
    .io_interrupt(LevelGateway_43_1_io_interrupt),
    .io_plic_valid(LevelGateway_43_1_io_plic_valid),
    .io_plic_ready(LevelGateway_43_1_io_plic_ready),
    .io_plic_complete(LevelGateway_43_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_44_1 (
    .clock(LevelGateway_44_1_clock),
    .reset(LevelGateway_44_1_reset),
    .io_interrupt(LevelGateway_44_1_io_interrupt),
    .io_plic_valid(LevelGateway_44_1_io_plic_valid),
    .io_plic_ready(LevelGateway_44_1_io_plic_ready),
    .io_plic_complete(LevelGateway_44_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_45_1 (
    .clock(LevelGateway_45_1_clock),
    .reset(LevelGateway_45_1_reset),
    .io_interrupt(LevelGateway_45_1_io_interrupt),
    .io_plic_valid(LevelGateway_45_1_io_plic_valid),
    .io_plic_ready(LevelGateway_45_1_io_plic_ready),
    .io_plic_complete(LevelGateway_45_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_46_1 (
    .clock(LevelGateway_46_1_clock),
    .reset(LevelGateway_46_1_reset),
    .io_interrupt(LevelGateway_46_1_io_interrupt),
    .io_plic_valid(LevelGateway_46_1_io_plic_valid),
    .io_plic_ready(LevelGateway_46_1_io_plic_ready),
    .io_plic_complete(LevelGateway_46_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_47_1 (
    .clock(LevelGateway_47_1_clock),
    .reset(LevelGateway_47_1_reset),
    .io_interrupt(LevelGateway_47_1_io_interrupt),
    .io_plic_valid(LevelGateway_47_1_io_plic_valid),
    .io_plic_ready(LevelGateway_47_1_io_plic_ready),
    .io_plic_complete(LevelGateway_47_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_48_1 (
    .clock(LevelGateway_48_1_clock),
    .reset(LevelGateway_48_1_reset),
    .io_interrupt(LevelGateway_48_1_io_interrupt),
    .io_plic_valid(LevelGateway_48_1_io_plic_valid),
    .io_plic_ready(LevelGateway_48_1_io_plic_ready),
    .io_plic_complete(LevelGateway_48_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_49_1 (
    .clock(LevelGateway_49_1_clock),
    .reset(LevelGateway_49_1_reset),
    .io_interrupt(LevelGateway_49_1_io_interrupt),
    .io_plic_valid(LevelGateway_49_1_io_plic_valid),
    .io_plic_ready(LevelGateway_49_1_io_plic_ready),
    .io_plic_complete(LevelGateway_49_1_io_plic_complete)
  );
  sirv_LevelGateway u_LevelGateway_50_1 (
    .clock(LevelGateway_50_1_clock),
    .reset(LevelGateway_50_1_reset),
    .io_interrupt(LevelGateway_50_1_io_interrupt),
    .io_plic_valid(LevelGateway_50_1_io_plic_valid),
    .io_plic_ready(LevelGateway_50_1_io_plic_ready),
    .io_plic_complete(LevelGateway_50_1_io_plic_complete)
  );
  assign io_tl_in_0_a_ready = T_3130_ready;
  assign io_tl_in_0_b_valid = 1'h0;
  assign io_tl_in_0_b_bits_opcode = GEN_60;
  assign io_tl_in_0_b_bits_param = GEN_91;
  assign io_tl_in_0_b_bits_size = GEN_143;
  assign io_tl_in_0_b_bits_source = GEN_364;
  assign io_tl_in_0_b_bits_address = GEN_3714;
  assign io_tl_in_0_b_bits_mask = GEN_3715;
  assign io_tl_in_0_b_bits_data = GEN_3716;
  assign io_tl_in_0_c_ready = 1'h1;
  assign io_tl_in_0_d_valid = T_3169_valid;
  assign io_tl_in_0_d_bits_opcode = {{2'd0}, T_3169_bits_read};
  assign io_tl_in_0_d_bits_param = T_49219_param;
  assign io_tl_in_0_d_bits_size = T_49219_size;
  assign io_tl_in_0_d_bits_source = T_49219_source;
  assign io_tl_in_0_d_bits_sink = T_49219_sink;
  assign io_tl_in_0_d_bits_addr_lo = T_49219_addr_lo;
  assign io_tl_in_0_d_bits_data = T_3169_bits_data;
  assign io_tl_in_0_d_bits_error = T_49219_error;
  assign io_tl_in_0_e_ready = 1'h1;
  assign io_harts_0_0 = T_3106;
  assign LevelGateway_51_clock = clock;
  assign LevelGateway_51_reset = reset;
  assign LevelGateway_51_io_interrupt = io_devices_0_0;
  assign LevelGateway_51_io_plic_ready = gateways_0_ready;
  assign LevelGateway_51_io_plic_complete = gateways_0_complete;
  assign LevelGateway_1_1_clock = clock;
  assign LevelGateway_1_1_reset = reset;
  assign LevelGateway_1_1_io_interrupt = io_devices_0_1;
  assign LevelGateway_1_1_io_plic_ready = gateways_1_ready;
  assign LevelGateway_1_1_io_plic_complete = gateways_1_complete;
  assign LevelGateway_2_1_clock = clock;
  assign LevelGateway_2_1_reset = reset;
  assign LevelGateway_2_1_io_interrupt = io_devices_0_2;
  assign LevelGateway_2_1_io_plic_ready = gateways_2_ready;
  assign LevelGateway_2_1_io_plic_complete = gateways_2_complete;
  assign LevelGateway_3_1_clock = clock;
  assign LevelGateway_3_1_reset = reset;
  assign LevelGateway_3_1_io_interrupt = io_devices_0_3;
  assign LevelGateway_3_1_io_plic_ready = gateways_3_ready;
  assign LevelGateway_3_1_io_plic_complete = gateways_3_complete;
  assign LevelGateway_4_1_clock = clock;
  assign LevelGateway_4_1_reset = reset;
  assign LevelGateway_4_1_io_interrupt = io_devices_0_4;
  assign LevelGateway_4_1_io_plic_ready = gateways_4_ready;
  assign LevelGateway_4_1_io_plic_complete = gateways_4_complete;
  assign LevelGateway_5_1_clock = clock;
  assign LevelGateway_5_1_reset = reset;
  assign LevelGateway_5_1_io_interrupt = io_devices_0_5;
  assign LevelGateway_5_1_io_plic_ready = gateways_5_ready;
  assign LevelGateway_5_1_io_plic_complete = gateways_5_complete;
  assign LevelGateway_6_1_clock = clock;
  assign LevelGateway_6_1_reset = reset;
  assign LevelGateway_6_1_io_interrupt = io_devices_0_6;
  assign LevelGateway_6_1_io_plic_ready = gateways_6_ready;
  assign LevelGateway_6_1_io_plic_complete = gateways_6_complete;
  assign LevelGateway_7_1_clock = clock;
  assign LevelGateway_7_1_reset = reset;
  assign LevelGateway_7_1_io_interrupt = io_devices_0_7;
  assign LevelGateway_7_1_io_plic_ready = gateways_7_ready;
  assign LevelGateway_7_1_io_plic_complete = gateways_7_complete;
  assign LevelGateway_8_1_clock = clock;
  assign LevelGateway_8_1_reset = reset;
  assign LevelGateway_8_1_io_interrupt = io_devices_0_8;
  assign LevelGateway_8_1_io_plic_ready = gateways_8_ready;
  assign LevelGateway_8_1_io_plic_complete = gateways_8_complete;
  assign LevelGateway_9_1_clock = clock;
  assign LevelGateway_9_1_reset = reset;
  assign LevelGateway_9_1_io_interrupt = io_devices_0_9;
  assign LevelGateway_9_1_io_plic_ready = gateways_9_ready;
  assign LevelGateway_9_1_io_plic_complete = gateways_9_complete;
  assign LevelGateway_10_1_clock = clock;
  assign LevelGateway_10_1_reset = reset;
  assign LevelGateway_10_1_io_interrupt = io_devices_0_10;
  assign LevelGateway_10_1_io_plic_ready = gateways_10_ready;
  assign LevelGateway_10_1_io_plic_complete = gateways_10_complete;
  assign LevelGateway_11_1_clock = clock;
  assign LevelGateway_11_1_reset = reset;
  assign LevelGateway_11_1_io_interrupt = io_devices_0_11;
  assign LevelGateway_11_1_io_plic_ready = gateways_11_ready;
  assign LevelGateway_11_1_io_plic_complete = gateways_11_complete;
  assign LevelGateway_12_1_clock = clock;
  assign LevelGateway_12_1_reset = reset;
  assign LevelGateway_12_1_io_interrupt = io_devices_0_12;
  assign LevelGateway_12_1_io_plic_ready = gateways_12_ready;
  assign LevelGateway_12_1_io_plic_complete = gateways_12_complete;
  assign LevelGateway_13_1_clock = clock;
  assign LevelGateway_13_1_reset = reset;
  assign LevelGateway_13_1_io_interrupt = io_devices_0_13;
  assign LevelGateway_13_1_io_plic_ready = gateways_13_ready;
  assign LevelGateway_13_1_io_plic_complete = gateways_13_complete;
  assign LevelGateway_14_1_clock = clock;
  assign LevelGateway_14_1_reset = reset;
  assign LevelGateway_14_1_io_interrupt = io_devices_0_14;
  assign LevelGateway_14_1_io_plic_ready = gateways_14_ready;
  assign LevelGateway_14_1_io_plic_complete = gateways_14_complete;
  assign LevelGateway_15_1_clock = clock;
  assign LevelGateway_15_1_reset = reset;
  assign LevelGateway_15_1_io_interrupt = io_devices_0_15;
  assign LevelGateway_15_1_io_plic_ready = gateways_15_ready;
  assign LevelGateway_15_1_io_plic_complete = gateways_15_complete;
  assign LevelGateway_16_1_clock = clock;
  assign LevelGateway_16_1_reset = reset;
  assign LevelGateway_16_1_io_interrupt = io_devices_0_16;
  assign LevelGateway_16_1_io_plic_ready = gateways_16_ready;
  assign LevelGateway_16_1_io_plic_complete = gateways_16_complete;
  assign LevelGateway_17_1_clock = clock;
  assign LevelGateway_17_1_reset = reset;
  assign LevelGateway_17_1_io_interrupt = io_devices_0_17;
  assign LevelGateway_17_1_io_plic_ready = gateways_17_ready;
  assign LevelGateway_17_1_io_plic_complete = gateways_17_complete;
  assign LevelGateway_18_1_clock = clock;
  assign LevelGateway_18_1_reset = reset;
  assign LevelGateway_18_1_io_interrupt = io_devices_0_18;
  assign LevelGateway_18_1_io_plic_ready = gateways_18_ready;
  assign LevelGateway_18_1_io_plic_complete = gateways_18_complete;
  assign LevelGateway_19_1_clock = clock;
  assign LevelGateway_19_1_reset = reset;
  assign LevelGateway_19_1_io_interrupt = io_devices_0_19;
  assign LevelGateway_19_1_io_plic_ready = gateways_19_ready;
  assign LevelGateway_19_1_io_plic_complete = gateways_19_complete;
  assign LevelGateway_20_1_clock = clock;
  assign LevelGateway_20_1_reset = reset;
  assign LevelGateway_20_1_io_interrupt = io_devices_0_20;
  assign LevelGateway_20_1_io_plic_ready = gateways_20_ready;
  assign LevelGateway_20_1_io_plic_complete = gateways_20_complete;
  assign LevelGateway_21_1_clock = clock;
  assign LevelGateway_21_1_reset = reset;
  assign LevelGateway_21_1_io_interrupt = io_devices_0_21;
  assign LevelGateway_21_1_io_plic_ready = gateways_21_ready;
  assign LevelGateway_21_1_io_plic_complete = gateways_21_complete;
  assign LevelGateway_22_1_clock = clock;
  assign LevelGateway_22_1_reset = reset;
  assign LevelGateway_22_1_io_interrupt = io_devices_0_22;
  assign LevelGateway_22_1_io_plic_ready = gateways_22_ready;
  assign LevelGateway_22_1_io_plic_complete = gateways_22_complete;
  assign LevelGateway_23_1_clock = clock;
  assign LevelGateway_23_1_reset = reset;
  assign LevelGateway_23_1_io_interrupt = io_devices_0_23;
  assign LevelGateway_23_1_io_plic_ready = gateways_23_ready;
  assign LevelGateway_23_1_io_plic_complete = gateways_23_complete;
  assign LevelGateway_24_1_clock = clock;
  assign LevelGateway_24_1_reset = reset;
  assign LevelGateway_24_1_io_interrupt = io_devices_0_24;
  assign LevelGateway_24_1_io_plic_ready = gateways_24_ready;
  assign LevelGateway_24_1_io_plic_complete = gateways_24_complete;
  assign LevelGateway_25_1_clock = clock;
  assign LevelGateway_25_1_reset = reset;
  assign LevelGateway_25_1_io_interrupt = io_devices_0_25;
  assign LevelGateway_25_1_io_plic_ready = gateways_25_ready;
  assign LevelGateway_25_1_io_plic_complete = gateways_25_complete;
  assign LevelGateway_26_1_clock = clock;
  assign LevelGateway_26_1_reset = reset;
  assign LevelGateway_26_1_io_interrupt = io_devices_0_26;
  assign LevelGateway_26_1_io_plic_ready = gateways_26_ready;
  assign LevelGateway_26_1_io_plic_complete = gateways_26_complete;
  assign LevelGateway_27_1_clock = clock;
  assign LevelGateway_27_1_reset = reset;
  assign LevelGateway_27_1_io_interrupt = io_devices_0_27;
  assign LevelGateway_27_1_io_plic_ready = gateways_27_ready;
  assign LevelGateway_27_1_io_plic_complete = gateways_27_complete;
  assign LevelGateway_28_1_clock = clock;
  assign LevelGateway_28_1_reset = reset;
  assign LevelGateway_28_1_io_interrupt = io_devices_0_28;
  assign LevelGateway_28_1_io_plic_ready = gateways_28_ready;
  assign LevelGateway_28_1_io_plic_complete = gateways_28_complete;
  assign LevelGateway_29_1_clock = clock;
  assign LevelGateway_29_1_reset = reset;
  assign LevelGateway_29_1_io_interrupt = io_devices_0_29;
  assign LevelGateway_29_1_io_plic_ready = gateways_29_ready;
  assign LevelGateway_29_1_io_plic_complete = gateways_29_complete;
  assign LevelGateway_30_1_clock = clock;
  assign LevelGateway_30_1_reset = reset;
  assign LevelGateway_30_1_io_interrupt = io_devices_0_30;
  assign LevelGateway_30_1_io_plic_ready = gateways_30_ready;
  assign LevelGateway_30_1_io_plic_complete = gateways_30_complete;
  assign LevelGateway_31_1_clock = clock;
  assign LevelGateway_31_1_reset = reset;
  assign LevelGateway_31_1_io_interrupt = io_devices_0_31;
  assign LevelGateway_31_1_io_plic_ready = gateways_31_ready;
  assign LevelGateway_31_1_io_plic_complete = gateways_31_complete;
  assign LevelGateway_32_1_clock = clock;
  assign LevelGateway_32_1_reset = reset;
  assign LevelGateway_32_1_io_interrupt = io_devices_0_32;
  assign LevelGateway_32_1_io_plic_ready = gateways_32_ready;
  assign LevelGateway_32_1_io_plic_complete = gateways_32_complete;
  assign LevelGateway_33_1_clock = clock;
  assign LevelGateway_33_1_reset = reset;
  assign LevelGateway_33_1_io_interrupt = io_devices_0_33;
  assign LevelGateway_33_1_io_plic_ready = gateways_33_ready;
  assign LevelGateway_33_1_io_plic_complete = gateways_33_complete;
  assign LevelGateway_34_1_clock = clock;
  assign LevelGateway_34_1_reset = reset;
  assign LevelGateway_34_1_io_interrupt = io_devices_0_34;
  assign LevelGateway_34_1_io_plic_ready = gateways_34_ready;
  assign LevelGateway_34_1_io_plic_complete = gateways_34_complete;
  assign LevelGateway_35_1_clock = clock;
  assign LevelGateway_35_1_reset = reset;
  assign LevelGateway_35_1_io_interrupt = io_devices_0_35;
  assign LevelGateway_35_1_io_plic_ready = gateways_35_ready;
  assign LevelGateway_35_1_io_plic_complete = gateways_35_complete;
  assign LevelGateway_36_1_clock = clock;
  assign LevelGateway_36_1_reset = reset;
  assign LevelGateway_36_1_io_interrupt = io_devices_0_36;
  assign LevelGateway_36_1_io_plic_ready = gateways_36_ready;
  assign LevelGateway_36_1_io_plic_complete = gateways_36_complete;
  assign LevelGateway_37_1_clock = clock;
  assign LevelGateway_37_1_reset = reset;
  assign LevelGateway_37_1_io_interrupt = io_devices_0_37;
  assign LevelGateway_37_1_io_plic_ready = gateways_37_ready;
  assign LevelGateway_37_1_io_plic_complete = gateways_37_complete;
  assign LevelGateway_38_1_clock = clock;
  assign LevelGateway_38_1_reset = reset;
  assign LevelGateway_38_1_io_interrupt = io_devices_0_38;
  assign LevelGateway_38_1_io_plic_ready = gateways_38_ready;
  assign LevelGateway_38_1_io_plic_complete = gateways_38_complete;
  assign LevelGateway_39_1_clock = clock;
  assign LevelGateway_39_1_reset = reset;
  assign LevelGateway_39_1_io_interrupt = io_devices_0_39;
  assign LevelGateway_39_1_io_plic_ready = gateways_39_ready;
  assign LevelGateway_39_1_io_plic_complete = gateways_39_complete;
  assign LevelGateway_40_1_clock = clock;
  assign LevelGateway_40_1_reset = reset;
  assign LevelGateway_40_1_io_interrupt = io_devices_0_40;
  assign LevelGateway_40_1_io_plic_ready = gateways_40_ready;
  assign LevelGateway_40_1_io_plic_complete = gateways_40_complete;
  assign LevelGateway_41_1_clock = clock;
  assign LevelGateway_41_1_reset = reset;
  assign LevelGateway_41_1_io_interrupt = io_devices_0_41;
  assign LevelGateway_41_1_io_plic_ready = gateways_41_ready;
  assign LevelGateway_41_1_io_plic_complete = gateways_41_complete;
  assign LevelGateway_42_1_clock = clock;
  assign LevelGateway_42_1_reset = reset;
  assign LevelGateway_42_1_io_interrupt = io_devices_0_42;
  assign LevelGateway_42_1_io_plic_ready = gateways_42_ready;
  assign LevelGateway_42_1_io_plic_complete = gateways_42_complete;
  assign LevelGateway_43_1_clock = clock;
  assign LevelGateway_43_1_reset = reset;
  assign LevelGateway_43_1_io_interrupt = io_devices_0_43;
  assign LevelGateway_43_1_io_plic_ready = gateways_43_ready;
  assign LevelGateway_43_1_io_plic_complete = gateways_43_complete;
  assign LevelGateway_44_1_clock = clock;
  assign LevelGateway_44_1_reset = reset;
  assign LevelGateway_44_1_io_interrupt = io_devices_0_44;
  assign LevelGateway_44_1_io_plic_ready = gateways_44_ready;
  assign LevelGateway_44_1_io_plic_complete = gateways_44_complete;
  assign LevelGateway_45_1_clock = clock;
  assign LevelGateway_45_1_reset = reset;
  assign LevelGateway_45_1_io_interrupt = io_devices_0_45;
  assign LevelGateway_45_1_io_plic_ready = gateways_45_ready;
  assign LevelGateway_45_1_io_plic_complete = gateways_45_complete;
  assign LevelGateway_46_1_clock = clock;
  assign LevelGateway_46_1_reset = reset;
  assign LevelGateway_46_1_io_interrupt = io_devices_0_46;
  assign LevelGateway_46_1_io_plic_ready = gateways_46_ready;
  assign LevelGateway_46_1_io_plic_complete = gateways_46_complete;
  assign LevelGateway_47_1_clock = clock;
  assign LevelGateway_47_1_reset = reset;
  assign LevelGateway_47_1_io_interrupt = io_devices_0_47;
  assign LevelGateway_47_1_io_plic_ready = gateways_47_ready;
  assign LevelGateway_47_1_io_plic_complete = gateways_47_complete;
  assign LevelGateway_48_1_clock = clock;
  assign LevelGateway_48_1_reset = reset;
  assign LevelGateway_48_1_io_interrupt = io_devices_0_48;
  assign LevelGateway_48_1_io_plic_ready = gateways_48_ready;
  assign LevelGateway_48_1_io_plic_complete = gateways_48_complete;
  assign LevelGateway_49_1_clock = clock;
  assign LevelGateway_49_1_reset = reset;
  assign LevelGateway_49_1_io_interrupt = io_devices_0_49;
  assign LevelGateway_49_1_io_plic_ready = gateways_49_ready;
  assign LevelGateway_49_1_io_plic_complete = gateways_49_complete;
  assign LevelGateway_50_1_clock = clock;
  assign LevelGateway_50_1_reset = reset;
  assign LevelGateway_50_1_io_interrupt = io_devices_0_50;
  assign LevelGateway_50_1_io_plic_ready = gateways_50_ready;
  assign LevelGateway_50_1_io_plic_complete = gateways_50_complete;
  assign gateways_0_valid = LevelGateway_51_io_plic_valid;
  assign gateways_0_ready = T_2485;
  assign gateways_0_complete = GEN_298;
  assign gateways_1_valid = LevelGateway_1_1_io_plic_valid;
  assign gateways_1_ready = T_2489;
  assign gateways_1_complete = GEN_299;
  assign gateways_2_valid = LevelGateway_2_1_io_plic_valid;
  assign gateways_2_ready = T_2493;
  assign gateways_2_complete = GEN_300;
  assign gateways_3_valid = LevelGateway_3_1_io_plic_valid;
  assign gateways_3_ready = T_2497;
  assign gateways_3_complete = GEN_301;
  assign gateways_4_valid = LevelGateway_4_1_io_plic_valid;
  assign gateways_4_ready = T_2501;
  assign gateways_4_complete = GEN_302;
  assign gateways_5_valid = LevelGateway_5_1_io_plic_valid;
  assign gateways_5_ready = T_2505;
  assign gateways_5_complete = GEN_303;
  assign gateways_6_valid = LevelGateway_6_1_io_plic_valid;
  assign gateways_6_ready = T_2509;
  assign gateways_6_complete = GEN_304;
  assign gateways_7_valid = LevelGateway_7_1_io_plic_valid;
  assign gateways_7_ready = T_2513;
  assign gateways_7_complete = GEN_305;
  assign gateways_8_valid = LevelGateway_8_1_io_plic_valid;
  assign gateways_8_ready = T_2517;
  assign gateways_8_complete = GEN_306;
  assign gateways_9_valid = LevelGateway_9_1_io_plic_valid;
  assign gateways_9_ready = T_2521;
  assign gateways_9_complete = GEN_307;
  assign gateways_10_valid = LevelGateway_10_1_io_plic_valid;
  assign gateways_10_ready = T_2525;
  assign gateways_10_complete = GEN_308;
  assign gateways_11_valid = LevelGateway_11_1_io_plic_valid;
  assign gateways_11_ready = T_2529;
  assign gateways_11_complete = GEN_309;
  assign gateways_12_valid = LevelGateway_12_1_io_plic_valid;
  assign gateways_12_ready = T_2533;
  assign gateways_12_complete = GEN_310;
  assign gateways_13_valid = LevelGateway_13_1_io_plic_valid;
  assign gateways_13_ready = T_2537;
  assign gateways_13_complete = GEN_311;
  assign gateways_14_valid = LevelGateway_14_1_io_plic_valid;
  assign gateways_14_ready = T_2541;
  assign gateways_14_complete = GEN_312;
  assign gateways_15_valid = LevelGateway_15_1_io_plic_valid;
  assign gateways_15_ready = T_2545;
  assign gateways_15_complete = GEN_313;
  assign gateways_16_valid = LevelGateway_16_1_io_plic_valid;
  assign gateways_16_ready = T_2549;
  assign gateways_16_complete = GEN_314;
  assign gateways_17_valid = LevelGateway_17_1_io_plic_valid;
  assign gateways_17_ready = T_2553;
  assign gateways_17_complete = GEN_315;
  assign gateways_18_valid = LevelGateway_18_1_io_plic_valid;
  assign gateways_18_ready = T_2557;
  assign gateways_18_complete = GEN_316;
  assign gateways_19_valid = LevelGateway_19_1_io_plic_valid;
  assign gateways_19_ready = T_2561;
  assign gateways_19_complete = GEN_317;
  assign gateways_20_valid = LevelGateway_20_1_io_plic_valid;
  assign gateways_20_ready = T_2565;
  assign gateways_20_complete = GEN_318;
  assign gateways_21_valid = LevelGateway_21_1_io_plic_valid;
  assign gateways_21_ready = T_2569;
  assign gateways_21_complete = GEN_319;
  assign gateways_22_valid = LevelGateway_22_1_io_plic_valid;
  assign gateways_22_ready = T_2573;
  assign gateways_22_complete = GEN_320;
  assign gateways_23_valid = LevelGateway_23_1_io_plic_valid;
  assign gateways_23_ready = T_2577;
  assign gateways_23_complete = GEN_321;
  assign gateways_24_valid = LevelGateway_24_1_io_plic_valid;
  assign gateways_24_ready = T_2581;
  assign gateways_24_complete = GEN_322;
  assign gateways_25_valid = LevelGateway_25_1_io_plic_valid;
  assign gateways_25_ready = T_2585;
  assign gateways_25_complete = GEN_323;
  assign gateways_26_valid = LevelGateway_26_1_io_plic_valid;
  assign gateways_26_ready = T_2589;
  assign gateways_26_complete = GEN_324;
  assign gateways_27_valid = LevelGateway_27_1_io_plic_valid;
  assign gateways_27_ready = T_2593;
  assign gateways_27_complete = GEN_325;
  assign gateways_28_valid = LevelGateway_28_1_io_plic_valid;
  assign gateways_28_ready = T_2597;
  assign gateways_28_complete = GEN_326;
  assign gateways_29_valid = LevelGateway_29_1_io_plic_valid;
  assign gateways_29_ready = T_2601;
  assign gateways_29_complete = GEN_327;
  assign gateways_30_valid = LevelGateway_30_1_io_plic_valid;
  assign gateways_30_ready = T_2605;
  assign gateways_30_complete = GEN_328;
  assign gateways_31_valid = LevelGateway_31_1_io_plic_valid;
  assign gateways_31_ready = T_2609;
  assign gateways_31_complete = GEN_329;
  assign gateways_32_valid = LevelGateway_32_1_io_plic_valid;
  assign gateways_32_ready = T_2613;
  assign gateways_32_complete = GEN_330;
  assign gateways_33_valid = LevelGateway_33_1_io_plic_valid;
  assign gateways_33_ready = T_2617;
  assign gateways_33_complete = GEN_331;
  assign gateways_34_valid = LevelGateway_34_1_io_plic_valid;
  assign gateways_34_ready = T_2621;
  assign gateways_34_complete = GEN_332;
  assign gateways_35_valid = LevelGateway_35_1_io_plic_valid;
  assign gateways_35_ready = T_2625;
  assign gateways_35_complete = GEN_333;
  assign gateways_36_valid = LevelGateway_36_1_io_plic_valid;
  assign gateways_36_ready = T_2629;
  assign gateways_36_complete = GEN_334;
  assign gateways_37_valid = LevelGateway_37_1_io_plic_valid;
  assign gateways_37_ready = T_2633;
  assign gateways_37_complete = GEN_335;
  assign gateways_38_valid = LevelGateway_38_1_io_plic_valid;
  assign gateways_38_ready = T_2637;
  assign gateways_38_complete = GEN_336;
  assign gateways_39_valid = LevelGateway_39_1_io_plic_valid;
  assign gateways_39_ready = T_2641;
  assign gateways_39_complete = GEN_337;
  assign gateways_40_valid = LevelGateway_40_1_io_plic_valid;
  assign gateways_40_ready = T_2645;
  assign gateways_40_complete = GEN_338;
  assign gateways_41_valid = LevelGateway_41_1_io_plic_valid;
  assign gateways_41_ready = T_2649;
  assign gateways_41_complete = GEN_339;
  assign gateways_42_valid = LevelGateway_42_1_io_plic_valid;
  assign gateways_42_ready = T_2653;
  assign gateways_42_complete = GEN_340;
  assign gateways_43_valid = LevelGateway_43_1_io_plic_valid;
  assign gateways_43_ready = T_2657;
  assign gateways_43_complete = GEN_341;
  assign gateways_44_valid = LevelGateway_44_1_io_plic_valid;
  assign gateways_44_ready = T_2661;
  assign gateways_44_complete = GEN_342;
  assign gateways_45_valid = LevelGateway_45_1_io_plic_valid;
  assign gateways_45_ready = T_2665;
  assign gateways_45_complete = GEN_343;
  assign gateways_46_valid = LevelGateway_46_1_io_plic_valid;
  assign gateways_46_ready = T_2669;
  assign gateways_46_complete = GEN_344;
  assign gateways_47_valid = LevelGateway_47_1_io_plic_valid;
  assign gateways_47_ready = T_2673;
  assign gateways_47_complete = GEN_345;
  assign gateways_48_valid = LevelGateway_48_1_io_plic_valid;
  assign gateways_48_ready = T_2677;
  assign gateways_48_complete = GEN_346;
  assign gateways_49_valid = LevelGateway_49_1_io_plic_valid;
  assign gateways_49_ready = T_2681;
  assign gateways_49_complete = GEN_347;
  assign gateways_50_valid = LevelGateway_50_1_io_plic_valid;
  assign gateways_50_ready = T_2685;
  assign gateways_50_complete = GEN_348;
  assign T_2365_0 = 1'h0;
  assign T_2365_1 = 1'h0;
  assign T_2365_2 = 1'h0;
  assign T_2365_3 = 1'h0;
  assign T_2365_4 = 1'h0;
  assign T_2365_5 = 1'h0;
  assign T_2365_6 = 1'h0;
  assign T_2365_7 = 1'h0;
  assign T_2365_8 = 1'h0;
  assign T_2365_9 = 1'h0;
  assign T_2365_10 = 1'h0;
  assign T_2365_11 = 1'h0;
  assign T_2365_12 = 1'h0;
  assign T_2365_13 = 1'h0;
  assign T_2365_14 = 1'h0;
  assign T_2365_15 = 1'h0;
  assign T_2365_16 = 1'h0;
  assign T_2365_17 = 1'h0;
  assign T_2365_18 = 1'h0;
  assign T_2365_19 = 1'h0;
  assign T_2365_20 = 1'h0;
  assign T_2365_21 = 1'h0;
  assign T_2365_22 = 1'h0;
  assign T_2365_23 = 1'h0;
  assign T_2365_24 = 1'h0;
  assign T_2365_25 = 1'h0;
  assign T_2365_26 = 1'h0;
  assign T_2365_27 = 1'h0;
  assign T_2365_28 = 1'h0;
  assign T_2365_29 = 1'h0;
  assign T_2365_30 = 1'h0;
  assign T_2365_31 = 1'h0;
  assign T_2365_32 = 1'h0;
  assign T_2365_33 = 1'h0;
  assign T_2365_34 = 1'h0;
  assign T_2365_35 = 1'h0;
  assign T_2365_36 = 1'h0;
  assign T_2365_37 = 1'h0;
  assign T_2365_38 = 1'h0;
  assign T_2365_39 = 1'h0;
  assign T_2365_40 = 1'h0;
  assign T_2365_41 = 1'h0;
  assign T_2365_42 = 1'h0;
  assign T_2365_43 = 1'h0;
  assign T_2365_44 = 1'h0;
  assign T_2365_45 = 1'h0;
  assign T_2365_46 = 1'h0;
  assign T_2365_47 = 1'h0;
  assign T_2365_48 = 1'h0;
  assign T_2365_49 = 1'h0;
  assign T_2365_50 = 1'h0;
  assign T_2365_51 = 1'h0;
  assign T_2485 = pending_1 == 1'h0;
  assign GEN_9 = gateways_0_valid ? 1'h1 : pending_1;
  assign T_2489 = pending_2 == 1'h0;
  assign GEN_10 = gateways_1_valid ? 1'h1 : pending_2;
  assign T_2493 = pending_3 == 1'h0;
  assign GEN_11 = gateways_2_valid ? 1'h1 : pending_3;
  assign T_2497 = pending_4 == 1'h0;
  assign GEN_12 = gateways_3_valid ? 1'h1 : pending_4;
  assign T_2501 = pending_5 == 1'h0;
  assign GEN_13 = gateways_4_valid ? 1'h1 : pending_5;
  assign T_2505 = pending_6 == 1'h0;
  assign GEN_14 = gateways_5_valid ? 1'h1 : pending_6;
  assign T_2509 = pending_7 == 1'h0;
  assign GEN_15 = gateways_6_valid ? 1'h1 : pending_7;
  assign T_2513 = pending_8 == 1'h0;
  assign GEN_16 = gateways_7_valid ? 1'h1 : pending_8;
  assign T_2517 = pending_9 == 1'h0;
  assign GEN_17 = gateways_8_valid ? 1'h1 : pending_9;
  assign T_2521 = pending_10 == 1'h0;
  assign GEN_18 = gateways_9_valid ? 1'h1 : pending_10;
  assign T_2525 = pending_11 == 1'h0;
  assign GEN_19 = gateways_10_valid ? 1'h1 : pending_11;
  assign T_2529 = pending_12 == 1'h0;
  assign GEN_20 = gateways_11_valid ? 1'h1 : pending_12;
  assign T_2533 = pending_13 == 1'h0;
  assign GEN_21 = gateways_12_valid ? 1'h1 : pending_13;
  assign T_2537 = pending_14 == 1'h0;
  assign GEN_22 = gateways_13_valid ? 1'h1 : pending_14;
  assign T_2541 = pending_15 == 1'h0;
  assign GEN_23 = gateways_14_valid ? 1'h1 : pending_15;
  assign T_2545 = pending_16 == 1'h0;
  assign GEN_24 = gateways_15_valid ? 1'h1 : pending_16;
  assign T_2549 = pending_17 == 1'h0;
  assign GEN_25 = gateways_16_valid ? 1'h1 : pending_17;
  assign T_2553 = pending_18 == 1'h0;
  assign GEN_26 = gateways_17_valid ? 1'h1 : pending_18;
  assign T_2557 = pending_19 == 1'h0;
  assign GEN_27 = gateways_18_valid ? 1'h1 : pending_19;
  assign T_2561 = pending_20 == 1'h0;
  assign GEN_28 = gateways_19_valid ? 1'h1 : pending_20;
  assign T_2565 = pending_21 == 1'h0;
  assign GEN_29 = gateways_20_valid ? 1'h1 : pending_21;
  assign T_2569 = pending_22 == 1'h0;
  assign GEN_30 = gateways_21_valid ? 1'h1 : pending_22;
  assign T_2573 = pending_23 == 1'h0;
  assign GEN_31 = gateways_22_valid ? 1'h1 : pending_23;
  assign T_2577 = pending_24 == 1'h0;
  assign GEN_32 = gateways_23_valid ? 1'h1 : pending_24;
  assign T_2581 = pending_25 == 1'h0;
  assign GEN_33 = gateways_24_valid ? 1'h1 : pending_25;
  assign T_2585 = pending_26 == 1'h0;
  assign GEN_34 = gateways_25_valid ? 1'h1 : pending_26;
  assign T_2589 = pending_27 == 1'h0;
  assign GEN_35 = gateways_26_valid ? 1'h1 : pending_27;
  assign T_2593 = pending_28 == 1'h0;
  assign GEN_36 = gateways_27_valid ? 1'h1 : pending_28;
  assign T_2597 = pending_29 == 1'h0;
  assign GEN_37 = gateways_28_valid ? 1'h1 : pending_29;
  assign T_2601 = pending_30 == 1'h0;
  assign GEN_38 = gateways_29_valid ? 1'h1 : pending_30;
  assign T_2605 = pending_31 == 1'h0;
  assign GEN_39 = gateways_30_valid ? 1'h1 : pending_31;
  assign T_2609 = pending_32 == 1'h0;
  assign GEN_40 = gateways_31_valid ? 1'h1 : pending_32;
  assign T_2613 = pending_33 == 1'h0;
  assign GEN_41 = gateways_32_valid ? 1'h1 : pending_33;
  assign T_2617 = pending_34 == 1'h0;
  assign GEN_42 = gateways_33_valid ? 1'h1 : pending_34;
  assign T_2621 = pending_35 == 1'h0;
  assign GEN_43 = gateways_34_valid ? 1'h1 : pending_35;
  assign T_2625 = pending_36 == 1'h0;
  assign GEN_44 = gateways_35_valid ? 1'h1 : pending_36;
  assign T_2629 = pending_37 == 1'h0;
  assign GEN_45 = gateways_36_valid ? 1'h1 : pending_37;
  assign T_2633 = pending_38 == 1'h0;
  assign GEN_46 = gateways_37_valid ? 1'h1 : pending_38;
  assign T_2637 = pending_39 == 1'h0;
  assign GEN_47 = gateways_38_valid ? 1'h1 : pending_39;
  assign T_2641 = pending_40 == 1'h0;
  assign GEN_48 = gateways_39_valid ? 1'h1 : pending_40;
  assign T_2645 = pending_41 == 1'h0;
  assign GEN_49 = gateways_40_valid ? 1'h1 : pending_41;
  assign T_2649 = pending_42 == 1'h0;
  assign GEN_50 = gateways_41_valid ? 1'h1 : pending_42;
  assign T_2653 = pending_43 == 1'h0;
  assign GEN_51 = gateways_42_valid ? 1'h1 : pending_43;
  assign T_2657 = pending_44 == 1'h0;
  assign GEN_52 = gateways_43_valid ? 1'h1 : pending_44;
  assign T_2661 = pending_45 == 1'h0;
  assign GEN_53 = gateways_44_valid ? 1'h1 : pending_45;
  assign T_2665 = pending_46 == 1'h0;
  assign GEN_54 = gateways_45_valid ? 1'h1 : pending_46;
  assign T_2669 = pending_47 == 1'h0;
  assign GEN_55 = gateways_46_valid ? 1'h1 : pending_47;
  assign T_2673 = pending_48 == 1'h0;
  assign GEN_56 = gateways_47_valid ? 1'h1 : pending_48;
  assign T_2677 = pending_49 == 1'h0;
  assign GEN_57 = gateways_48_valid ? 1'h1 : pending_49;
  assign T_2681 = pending_50 == 1'h0;
  assign GEN_58 = gateways_49_valid ? 1'h1 : pending_50;
  assign T_2685 = pending_51 == 1'h0;
  assign GEN_59 = gateways_50_valid ? 1'h1 : pending_51;
  assign T_2692 = pending_1 & enables_0_1;
  assign T_2693 = {T_2692,priority_1};
  assign T_2694 = pending_2 & enables_0_2;
  assign T_2695 = {T_2694,priority_2};
  assign T_2696 = pending_3 & enables_0_3;
  assign T_2697 = {T_2696,priority_3};
  assign T_2698 = pending_4 & enables_0_4;
  assign T_2699 = {T_2698,priority_4};
  assign T_2700 = pending_5 & enables_0_5;
  assign T_2701 = {T_2700,priority_5};
  assign T_2702 = pending_6 & enables_0_6;
  assign T_2703 = {T_2702,priority_6};
  assign T_2704 = pending_7 & enables_0_7;
  assign T_2705 = {T_2704,priority_7};
  assign T_2706 = pending_8 & enables_0_8;
  assign T_2707 = {T_2706,priority_8};
  assign T_2708 = pending_9 & enables_0_9;
  assign T_2709 = {T_2708,priority_9};
  assign T_2710 = pending_10 & enables_0_10;
  assign T_2711 = {T_2710,priority_10};
  assign T_2712 = pending_11 & enables_0_11;
  assign T_2713 = {T_2712,priority_11};
  assign T_2714 = pending_12 & enables_0_12;
  assign T_2715 = {T_2714,priority_12};
  assign T_2716 = pending_13 & enables_0_13;
  assign T_2717 = {T_2716,priority_13};
  assign T_2718 = pending_14 & enables_0_14;
  assign T_2719 = {T_2718,priority_14};
  assign T_2720 = pending_15 & enables_0_15;
  assign T_2721 = {T_2720,priority_15};
  assign T_2722 = pending_16 & enables_0_16;
  assign T_2723 = {T_2722,priority_16};
  assign T_2724 = pending_17 & enables_0_17;
  assign T_2725 = {T_2724,priority_17};
  assign T_2726 = pending_18 & enables_0_18;
  assign T_2727 = {T_2726,priority_18};
  assign T_2728 = pending_19 & enables_0_19;
  assign T_2729 = {T_2728,priority_19};
  assign T_2730 = pending_20 & enables_0_20;
  assign T_2731 = {T_2730,priority_20};
  assign T_2732 = pending_21 & enables_0_21;
  assign T_2733 = {T_2732,priority_21};
  assign T_2734 = pending_22 & enables_0_22;
  assign T_2735 = {T_2734,priority_22};
  assign T_2736 = pending_23 & enables_0_23;
  assign T_2737 = {T_2736,priority_23};
  assign T_2738 = pending_24 & enables_0_24;
  assign T_2739 = {T_2738,priority_24};
  assign T_2740 = pending_25 & enables_0_25;
  assign T_2741 = {T_2740,priority_25};
  assign T_2742 = pending_26 & enables_0_26;
  assign T_2743 = {T_2742,priority_26};
  assign T_2744 = pending_27 & enables_0_27;
  assign T_2745 = {T_2744,priority_27};
  assign T_2746 = pending_28 & enables_0_28;
  assign T_2747 = {T_2746,priority_28};
  assign T_2748 = pending_29 & enables_0_29;
  assign T_2749 = {T_2748,priority_29};
  assign T_2750 = pending_30 & enables_0_30;
  assign T_2751 = {T_2750,priority_30};
  assign T_2752 = pending_31 & enables_0_31;
  assign T_2753 = {T_2752,priority_31};
  assign T_2754 = pending_32 & enables_0_32;
  assign T_2755 = {T_2754,priority_32};
  assign T_2756 = pending_33 & enables_0_33;
  assign T_2757 = {T_2756,priority_33};
  assign T_2758 = pending_34 & enables_0_34;
  assign T_2759 = {T_2758,priority_34};
  assign T_2760 = pending_35 & enables_0_35;
  assign T_2761 = {T_2760,priority_35};
  assign T_2762 = pending_36 & enables_0_36;
  assign T_2763 = {T_2762,priority_36};
  assign T_2764 = pending_37 & enables_0_37;
  assign T_2765 = {T_2764,priority_37};
  assign T_2766 = pending_38 & enables_0_38;
  assign T_2767 = {T_2766,priority_38};
  assign T_2768 = pending_39 & enables_0_39;
  assign T_2769 = {T_2768,priority_39};
  assign T_2770 = pending_40 & enables_0_40;
  assign T_2771 = {T_2770,priority_40};
  assign T_2772 = pending_41 & enables_0_41;
  assign T_2773 = {T_2772,priority_41};
  assign T_2774 = pending_42 & enables_0_42;
  assign T_2775 = {T_2774,priority_42};
  assign T_2776 = pending_43 & enables_0_43;
  assign T_2777 = {T_2776,priority_43};
  assign T_2778 = pending_44 & enables_0_44;
  assign T_2779 = {T_2778,priority_44};
  assign T_2780 = pending_45 & enables_0_45;
  assign T_2781 = {T_2780,priority_45};
  assign T_2782 = pending_46 & enables_0_46;
  assign T_2783 = {T_2782,priority_46};
  assign T_2784 = pending_47 & enables_0_47;
  assign T_2785 = {T_2784,priority_47};
  assign T_2786 = pending_48 & enables_0_48;
  assign T_2787 = {T_2786,priority_48};
  assign T_2788 = pending_49 & enables_0_49;
  assign T_2789 = {T_2788,priority_49};
  assign T_2790 = pending_50 & enables_0_50;
  assign T_2791 = {T_2790,priority_50};
  assign T_2792 = pending_51 & enables_0_51;
  assign T_2793 = {T_2792,priority_51};
  assign T_2798 = 4'h8 >= T_2693;
  assign T_2799 = T_2798 ? 4'h8 : T_2693;
  assign T_2802 = T_2798 ? 1'h0 : 1'h1;
  assign T_2805 = T_2695 >= T_2697;
  assign T_2806 = T_2805 ? T_2695 : T_2697;
  assign T_2809 = T_2805 ? 1'h0 : 1'h1;
  assign T_2810 = T_2799 >= T_2806;
  assign T_2811 = T_2810 ? T_2799 : T_2806;
  assign GEN_3489 = {{1'd0}, T_2809};
  assign T_2813 = 2'h2 | GEN_3489;
  assign T_2814 = T_2810 ? {{1'd0}, T_2802} : T_2813;
  assign T_2817 = T_2699 >= T_2701;
  assign T_2818 = T_2817 ? T_2699 : T_2701;
  assign T_2821 = T_2817 ? 1'h0 : 1'h1;
  assign T_2824 = T_2703 >= T_2705;
  assign T_2825 = T_2824 ? T_2703 : T_2705;
  assign T_2828 = T_2824 ? 1'h0 : 1'h1;
  assign T_2829 = T_2818 >= T_2825;
  assign T_2830 = T_2829 ? T_2818 : T_2825;
  assign GEN_3490 = {{1'd0}, T_2828};
  assign T_2832 = 2'h2 | GEN_3490;
  assign T_2833 = T_2829 ? {{1'd0}, T_2821} : T_2832;
  assign T_2834 = T_2811 >= T_2830;
  assign T_2835 = T_2834 ? T_2811 : T_2830;
  assign GEN_3491 = {{1'd0}, T_2833};
  assign T_2837 = 3'h4 | GEN_3491;
  assign T_2838 = T_2834 ? {{1'd0}, T_2814} : T_2837;
  assign T_2841 = T_2707 >= T_2709;
  assign T_2842 = T_2841 ? T_2707 : T_2709;
  assign T_2845 = T_2841 ? 1'h0 : 1'h1;
  assign T_2848 = T_2711 >= T_2713;
  assign T_2849 = T_2848 ? T_2711 : T_2713;
  assign T_2852 = T_2848 ? 1'h0 : 1'h1;
  assign T_2853 = T_2842 >= T_2849;
  assign T_2854 = T_2853 ? T_2842 : T_2849;
  assign GEN_3492 = {{1'd0}, T_2852};
  assign T_2856 = 2'h2 | GEN_3492;
  assign T_2857 = T_2853 ? {{1'd0}, T_2845} : T_2856;
  assign T_2860 = T_2715 >= T_2717;
  assign T_2861 = T_2860 ? T_2715 : T_2717;
  assign T_2864 = T_2860 ? 1'h0 : 1'h1;
  assign T_2867 = T_2719 >= T_2721;
  assign T_2868 = T_2867 ? T_2719 : T_2721;
  assign T_2871 = T_2867 ? 1'h0 : 1'h1;
  assign T_2872 = T_2861 >= T_2868;
  assign T_2873 = T_2872 ? T_2861 : T_2868;
  assign GEN_3493 = {{1'd0}, T_2871};
  assign T_2875 = 2'h2 | GEN_3493;
  assign T_2876 = T_2872 ? {{1'd0}, T_2864} : T_2875;
  assign T_2877 = T_2854 >= T_2873;
  assign T_2878 = T_2877 ? T_2854 : T_2873;
  assign GEN_3494 = {{1'd0}, T_2876};
  assign T_2880 = 3'h4 | GEN_3494;
  assign T_2881 = T_2877 ? {{1'd0}, T_2857} : T_2880;
  assign T_2882 = T_2835 >= T_2878;
  assign T_2883 = T_2882 ? T_2835 : T_2878;
  assign GEN_3495 = {{1'd0}, T_2881};
  assign T_2885 = 4'h8 | GEN_3495;
  assign T_2886 = T_2882 ? {{1'd0}, T_2838} : T_2885;
  assign T_2889 = T_2723 >= T_2725;
  assign T_2890 = T_2889 ? T_2723 : T_2725;
  assign T_2893 = T_2889 ? 1'h0 : 1'h1;
  assign T_2896 = T_2727 >= T_2729;
  assign T_2897 = T_2896 ? T_2727 : T_2729;
  assign T_2900 = T_2896 ? 1'h0 : 1'h1;
  assign T_2901 = T_2890 >= T_2897;
  assign T_2902 = T_2901 ? T_2890 : T_2897;
  assign GEN_3496 = {{1'd0}, T_2900};
  assign T_2904 = 2'h2 | GEN_3496;
  assign T_2905 = T_2901 ? {{1'd0}, T_2893} : T_2904;
  assign T_2908 = T_2731 >= T_2733;
  assign T_2909 = T_2908 ? T_2731 : T_2733;
  assign T_2912 = T_2908 ? 1'h0 : 1'h1;
  assign T_2915 = T_2735 >= T_2737;
  assign T_2916 = T_2915 ? T_2735 : T_2737;
  assign T_2919 = T_2915 ? 1'h0 : 1'h1;
  assign T_2920 = T_2909 >= T_2916;
  assign T_2921 = T_2920 ? T_2909 : T_2916;
  assign GEN_3497 = {{1'd0}, T_2919};
  assign T_2923 = 2'h2 | GEN_3497;
  assign T_2924 = T_2920 ? {{1'd0}, T_2912} : T_2923;
  assign T_2925 = T_2902 >= T_2921;
  assign T_2926 = T_2925 ? T_2902 : T_2921;
  assign GEN_3498 = {{1'd0}, T_2924};
  assign T_2928 = 3'h4 | GEN_3498;
  assign T_2929 = T_2925 ? {{1'd0}, T_2905} : T_2928;
  assign T_2932 = T_2739 >= T_2741;
  assign T_2933 = T_2932 ? T_2739 : T_2741;
  assign T_2936 = T_2932 ? 1'h0 : 1'h1;
  assign T_2939 = T_2743 >= T_2745;
  assign T_2940 = T_2939 ? T_2743 : T_2745;
  assign T_2943 = T_2939 ? 1'h0 : 1'h1;
  assign T_2944 = T_2933 >= T_2940;
  assign T_2945 = T_2944 ? T_2933 : T_2940;
  assign GEN_3499 = {{1'd0}, T_2943};
  assign T_2947 = 2'h2 | GEN_3499;
  assign T_2948 = T_2944 ? {{1'd0}, T_2936} : T_2947;
  assign T_2951 = T_2747 >= T_2749;
  assign T_2952 = T_2951 ? T_2747 : T_2749;
  assign T_2955 = T_2951 ? 1'h0 : 1'h1;
  assign T_2958 = T_2751 >= T_2753;
  assign T_2959 = T_2958 ? T_2751 : T_2753;
  assign T_2962 = T_2958 ? 1'h0 : 1'h1;
  assign T_2963 = T_2952 >= T_2959;
  assign T_2964 = T_2963 ? T_2952 : T_2959;
  assign GEN_3500 = {{1'd0}, T_2962};
  assign T_2966 = 2'h2 | GEN_3500;
  assign T_2967 = T_2963 ? {{1'd0}, T_2955} : T_2966;
  assign T_2968 = T_2945 >= T_2964;
  assign T_2969 = T_2968 ? T_2945 : T_2964;
  assign GEN_3501 = {{1'd0}, T_2967};
  assign T_2971 = 3'h4 | GEN_3501;
  assign T_2972 = T_2968 ? {{1'd0}, T_2948} : T_2971;
  assign T_2973 = T_2926 >= T_2969;
  assign T_2974 = T_2973 ? T_2926 : T_2969;
  assign GEN_3502 = {{1'd0}, T_2972};
  assign T_2976 = 4'h8 | GEN_3502;
  assign T_2977 = T_2973 ? {{1'd0}, T_2929} : T_2976;
  assign T_2978 = T_2883 >= T_2974;
  assign T_2979 = T_2978 ? T_2883 : T_2974;
  assign GEN_3503 = {{1'd0}, T_2977};
  assign T_2981 = 5'h10 | GEN_3503;
  assign T_2982 = T_2978 ? {{1'd0}, T_2886} : T_2981;
  assign T_2985 = T_2755 >= T_2757;
  assign T_2986 = T_2985 ? T_2755 : T_2757;
  assign T_2989 = T_2985 ? 1'h0 : 1'h1;
  assign T_2992 = T_2759 >= T_2761;
  assign T_2993 = T_2992 ? T_2759 : T_2761;
  assign T_2996 = T_2992 ? 1'h0 : 1'h1;
  assign T_2997 = T_2986 >= T_2993;
  assign T_2998 = T_2997 ? T_2986 : T_2993;
  assign GEN_3504 = {{1'd0}, T_2996};
  assign T_3000 = 2'h2 | GEN_3504;
  assign T_3001 = T_2997 ? {{1'd0}, T_2989} : T_3000;
  assign T_3004 = T_2763 >= T_2765;
  assign T_3005 = T_3004 ? T_2763 : T_2765;
  assign T_3008 = T_3004 ? 1'h0 : 1'h1;
  assign T_3011 = T_2767 >= T_2769;
  assign T_3012 = T_3011 ? T_2767 : T_2769;
  assign T_3015 = T_3011 ? 1'h0 : 1'h1;
  assign T_3016 = T_3005 >= T_3012;
  assign T_3017 = T_3016 ? T_3005 : T_3012;
  assign GEN_3505 = {{1'd0}, T_3015};
  assign T_3019 = 2'h2 | GEN_3505;
  assign T_3020 = T_3016 ? {{1'd0}, T_3008} : T_3019;
  assign T_3021 = T_2998 >= T_3017;
  assign T_3022 = T_3021 ? T_2998 : T_3017;
  assign GEN_3506 = {{1'd0}, T_3020};
  assign T_3024 = 3'h4 | GEN_3506;
  assign T_3025 = T_3021 ? {{1'd0}, T_3001} : T_3024;
  assign T_3028 = T_2771 >= T_2773;
  assign T_3029 = T_3028 ? T_2771 : T_2773;
  assign T_3032 = T_3028 ? 1'h0 : 1'h1;
  assign T_3035 = T_2775 >= T_2777;
  assign T_3036 = T_3035 ? T_2775 : T_2777;
  assign T_3039 = T_3035 ? 1'h0 : 1'h1;
  assign T_3040 = T_3029 >= T_3036;
  assign T_3041 = T_3040 ? T_3029 : T_3036;
  assign GEN_3507 = {{1'd0}, T_3039};
  assign T_3043 = 2'h2 | GEN_3507;
  assign T_3044 = T_3040 ? {{1'd0}, T_3032} : T_3043;
  assign T_3047 = T_2779 >= T_2781;
  assign T_3048 = T_3047 ? T_2779 : T_2781;
  assign T_3051 = T_3047 ? 1'h0 : 1'h1;
  assign T_3054 = T_2783 >= T_2785;
  assign T_3055 = T_3054 ? T_2783 : T_2785;
  assign T_3058 = T_3054 ? 1'h0 : 1'h1;
  assign T_3059 = T_3048 >= T_3055;
  assign T_3060 = T_3059 ? T_3048 : T_3055;
  assign GEN_3508 = {{1'd0}, T_3058};
  assign T_3062 = 2'h2 | GEN_3508;
  assign T_3063 = T_3059 ? {{1'd0}, T_3051} : T_3062;
  assign T_3064 = T_3041 >= T_3060;
  assign T_3065 = T_3064 ? T_3041 : T_3060;
  assign GEN_3509 = {{1'd0}, T_3063};
  assign T_3067 = 3'h4 | GEN_3509;
  assign T_3068 = T_3064 ? {{1'd0}, T_3044} : T_3067;
  assign T_3069 = T_3022 >= T_3065;
  assign T_3070 = T_3069 ? T_3022 : T_3065;
  assign GEN_3510 = {{1'd0}, T_3068};
  assign T_3072 = 4'h8 | GEN_3510;
  assign T_3073 = T_3069 ? {{1'd0}, T_3025} : T_3072;
  assign T_3076 = T_2787 >= T_2789;
  assign T_3077 = T_3076 ? T_2787 : T_2789;
  assign T_3080 = T_3076 ? 1'h0 : 1'h1;
  assign T_3083 = T_2791 >= T_2793;
  assign T_3084 = T_3083 ? T_2791 : T_2793;
  assign T_3087 = T_3083 ? 1'h0 : 1'h1;
  assign T_3088 = T_3077 >= T_3084;
  assign T_3089 = T_3088 ? T_3077 : T_3084;
  assign GEN_3511 = {{1'd0}, T_3087};
  assign T_3091 = 2'h2 | GEN_3511;
  assign T_3092 = T_3088 ? {{1'd0}, T_3080} : T_3091;
  assign T_3093 = T_3070 >= T_3089;
  assign T_3094 = T_3093 ? T_3070 : T_3089;
  assign GEN_3512 = {{3'd0}, T_3092};
  assign T_3096 = 5'h10 | GEN_3512;
  assign T_3097 = T_3093 ? {{1'd0}, T_3073} : T_3096;
  assign T_3098 = T_2979 >= T_3094;
  assign T_3099 = T_3098 ? T_2979 : T_3094;
  assign GEN_3513 = {{1'd0}, T_3097};
  assign T_3101 = 6'h20 | GEN_3513;
  assign T_3102 = T_3098 ? {{1'd0}, T_2982} : T_3101;
  assign T_3105 = {1'h1,threshold_0};
  assign T_3106 = T_3103 > T_3105;
  assign T_3130_ready = T_24261;
  assign T_3130_valid = io_tl_in_0_a_valid;
  assign T_3130_bits_read = T_3147;
  assign T_3130_bits_index = T_3148[23:0];
  assign T_3130_bits_data = io_tl_in_0_a_bits_data;
  assign T_3130_bits_mask = io_tl_in_0_a_bits_mask;
  assign T_3130_bits_extra = T_3151;
  assign T_3147 = io_tl_in_0_a_bits_opcode == 3'h4;
  assign T_3148 = io_tl_in_0_a_bits_address[27:2];
  assign T_3149 = io_tl_in_0_a_bits_address[1:0];
  assign T_3150 = {T_3149,io_tl_in_0_a_bits_source};
  assign T_3151 = {T_3150,io_tl_in_0_a_bits_size};
  assign T_3169_ready = io_tl_in_0_d_ready;
  assign T_3169_valid = T_24264;
  assign T_3169_bits_read = T_3205_bits_read;
  assign T_3169_bits_data = T_49204;
  assign T_3169_bits_extra = T_3205_bits_extra;
  assign T_3205_ready = T_24263;
  assign T_3205_valid = T_24262;
  assign T_3205_bits_read = T_3130_bits_read;
  assign T_3205_bits_index = T_3130_bits_index;
  assign T_3205_bits_data = T_3130_bits_data;
  assign T_3205_bits_mask = T_3130_bits_mask;
  assign T_3205_bits_extra = T_3130_bits_extra;
  assign T_4309_0 = T_35563;
  assign T_4309_1 = T_35691;
  assign T_4309_2 = T_35819;
  assign T_4309_3 = T_35947;
  assign T_4309_4 = T_36075;
  assign T_4309_5 = T_36203;
  assign T_4309_6 = T_36331;
  assign T_4309_7 = T_36459;
  assign T_4309_8 = T_36587;
  assign T_4309_9 = T_36715;
  assign T_4309_10 = T_36843;
  assign T_4309_11 = T_36971;
  assign T_4309_12 = T_37099;
  assign T_4309_13 = T_37227;
  assign T_4309_14 = T_37355;
  assign T_4309_15 = T_37483;
  assign T_4309_16 = T_37611;
  assign T_4309_17 = T_37739;
  assign T_4309_18 = T_37867;
  assign T_4309_19 = T_37995;
  assign T_4309_20 = T_38123;
  assign T_4309_21 = T_38251;
  assign T_4309_22 = T_38379;
  assign T_4309_23 = T_38507;
  assign T_4309_24 = T_38635;
  assign T_4309_25 = T_38763;
  assign T_4309_26 = T_38891;
  assign T_4309_27 = T_39019;
  assign T_4309_28 = T_39147;
  assign T_4309_29 = T_39275;
  assign T_4309_30 = T_39403;
  assign T_4309_31 = T_39531;
  assign T_4309_32 = T_25296;
  assign T_4309_33 = T_25396;
  assign T_4309_34 = T_25496;
  assign T_4309_35 = T_26136;
  assign T_4309_36 = T_25776;
  assign T_4309_37 = T_26036;
  assign T_4309_38 = T_25796;
  assign T_4309_39 = T_25576;
  assign T_4309_40 = T_25696;
  assign T_4309_41 = T_39683;
  assign T_4309_42 = T_39763;
  assign T_4309_43 = T_39843;
  assign T_4309_44 = T_39923;
  assign T_4309_45 = T_40003;
  assign T_4309_46 = T_40083;
  assign T_4309_47 = T_40163;
  assign T_4309_48 = T_40243;
  assign T_4309_49 = T_40323;
  assign T_4309_50 = T_40403;
  assign T_4309_51 = T_40483;
  assign T_4309_52 = T_40563;
  assign T_4309_53 = T_40643;
  assign T_4309_54 = T_40723;
  assign T_4309_55 = T_40803;
  assign T_4309_56 = T_40883;
  assign T_4309_57 = T_40963;
  assign T_4309_58 = T_41043;
  assign T_4309_59 = T_41123;
  assign T_4309_60 = T_41203;
  assign T_4309_61 = T_26216;
  assign T_4309_62 = T_25876;
  assign T_4309_63 = T_30436;
  assign T_4309_64 = T_25316;
  assign T_4309_65 = T_25416;
  assign T_4309_66 = T_25856;
  assign T_4309_67 = T_26056;
  assign T_4309_68 = T_25716;
  assign T_4309_69 = T_25956;
  assign T_4309_70 = T_25476;
  assign T_4309_71 = T_25556;
  assign T_4309_72 = T_26116;
  assign T_4309_73 = T_25336;
  assign T_4309_74 = T_25936;
  assign T_4309_75 = T_25976;
  assign T_4309_76 = T_26196;
  assign T_4309_77 = T_25636;
  assign T_4309_78 = T_30416;
  assign T_4309_79 = T_41367;
  assign T_4309_80 = T_41495;
  assign T_4309_81 = T_41623;
  assign T_4309_82 = T_41751;
  assign T_4309_83 = T_41879;
  assign T_4309_84 = T_42007;
  assign T_4309_85 = T_42135;
  assign T_4309_86 = T_42263;
  assign T_4309_87 = T_42391;
  assign T_4309_88 = T_42519;
  assign T_4309_89 = T_42647;
  assign T_4309_90 = T_42775;
  assign T_4309_91 = T_42903;
  assign T_4309_92 = T_43031;
  assign T_4309_93 = T_43159;
  assign T_4309_94 = T_43287;
  assign T_4309_95 = T_43415;
  assign T_4309_96 = T_43543;
  assign T_4309_97 = T_43671;
  assign T_4309_98 = T_43799;
  assign T_4309_99 = T_43927;
  assign T_4309_100 = T_44055;
  assign T_4309_101 = T_44183;
  assign T_4309_102 = T_44311;
  assign T_4309_103 = T_44439;
  assign T_4309_104 = T_44567;
  assign T_4309_105 = T_44695;
  assign T_4309_106 = T_44823;
  assign T_4309_107 = T_44951;
  assign T_4309_108 = T_45079;
  assign T_4309_109 = T_45207;
  assign T_4309_110 = T_45335;
  assign T_4309_111 = T_25736;
  assign T_4309_112 = T_26176;
  assign T_4309_113 = T_25836;
  assign T_4309_114 = T_25536;
  assign T_4309_115 = T_26276;
  assign T_4309_116 = T_25436;
  assign T_4309_117 = T_26076;
  assign T_4309_118 = T_25356;
  assign T_4309_119 = T_25996;
  assign T_4309_120 = T_26256;
  assign T_4309_121 = T_45491;
  assign T_4309_122 = T_45571;
  assign T_4309_123 = T_45651;
  assign T_4309_124 = T_45731;
  assign T_4309_125 = T_45811;
  assign T_4309_126 = T_45891;
  assign T_4309_127 = T_45971;
  assign T_4309_128 = T_46051;
  assign T_4309_129 = T_46131;
  assign T_4309_130 = T_46211;
  assign T_4309_131 = T_46291;
  assign T_4309_132 = T_46371;
  assign T_4309_133 = T_46451;
  assign T_4309_134 = T_46531;
  assign T_4309_135 = T_46611;
  assign T_4309_136 = T_46691;
  assign T_4309_137 = T_46771;
  assign T_4309_138 = T_46851;
  assign T_4309_139 = T_46931;
  assign T_4309_140 = T_47011;
  assign T_4309_141 = T_25656;
  assign T_4309_142 = T_26296;
  assign T_4309_143 = T_25616;
  assign T_4309_144 = T_25916;
  assign T_4309_145 = T_25516;
  assign T_4309_146 = T_26156;
  assign T_4309_147 = T_26096;
  assign T_4309_148 = T_25816;
  assign T_4309_149 = T_25756;
  assign T_4309_150 = T_25456;
  assign T_4309_151 = T_26016;
  assign T_4309_152 = T_25896;
  assign T_4309_153 = T_26316;
  assign T_4309_154 = T_25676;
  assign T_4309_155 = T_25376;
  assign T_4309_156 = T_26236;
  assign T_4309_157 = T_25596;
  assign T_4314_0 = T_35595;
  assign T_4314_1 = T_35723;
  assign T_4314_2 = T_35851;
  assign T_4314_3 = T_35979;
  assign T_4314_4 = T_36107;
  assign T_4314_5 = T_36235;
  assign T_4314_6 = T_36363;
  assign T_4314_7 = T_36491;
  assign T_4314_8 = T_36619;
  assign T_4314_9 = T_36747;
  assign T_4314_10 = T_36875;
  assign T_4314_11 = T_37003;
  assign T_4314_12 = T_37131;
  assign T_4314_13 = T_37259;
  assign T_4314_14 = T_37387;
  assign T_4314_15 = T_37515;
  assign T_4314_16 = T_37643;
  assign T_4314_17 = T_37771;
  assign T_4314_18 = T_37899;
  assign T_4314_19 = T_38027;
  assign T_4314_20 = T_38155;
  assign T_4314_21 = T_38283;
  assign T_4314_22 = T_38411;
  assign T_4314_23 = T_38539;
  assign T_4314_24 = T_38667;
  assign T_4314_25 = T_38795;
  assign T_4314_26 = T_38923;
  assign T_4314_27 = T_39051;
  assign T_4314_28 = T_39179;
  assign T_4314_29 = T_39307;
  assign T_4314_30 = T_39435;
  assign T_4314_31 = T_39563;
  assign T_4314_32 = T_25302;
  assign T_4314_33 = T_25402;
  assign T_4314_34 = T_25502;
  assign T_4314_35 = T_26142;
  assign T_4314_36 = T_25782;
  assign T_4314_37 = T_26042;
  assign T_4314_38 = T_25802;
  assign T_4314_39 = T_25582;
  assign T_4314_40 = T_25702;
  assign T_4314_41 = T_39703;
  assign T_4314_42 = T_39783;
  assign T_4314_43 = T_39863;
  assign T_4314_44 = T_39943;
  assign T_4314_45 = T_40023;
  assign T_4314_46 = T_40103;
  assign T_4314_47 = T_40183;
  assign T_4314_48 = T_40263;
  assign T_4314_49 = T_40343;
  assign T_4314_50 = T_40423;
  assign T_4314_51 = T_40503;
  assign T_4314_52 = T_40583;
  assign T_4314_53 = T_40663;
  assign T_4314_54 = T_40743;
  assign T_4314_55 = T_40823;
  assign T_4314_56 = T_40903;
  assign T_4314_57 = T_40983;
  assign T_4314_58 = T_41063;
  assign T_4314_59 = T_41143;
  assign T_4314_60 = T_41223;
  assign T_4314_61 = T_26222;
  assign T_4314_62 = T_25882;
  assign T_4314_63 = T_30442;
  assign T_4314_64 = T_25322;
  assign T_4314_65 = T_25422;
  assign T_4314_66 = T_25862;
  assign T_4314_67 = T_26062;
  assign T_4314_68 = T_25722;
  assign T_4314_69 = T_25962;
  assign T_4314_70 = T_25482;
  assign T_4314_71 = T_25562;
  assign T_4314_72 = T_26122;
  assign T_4314_73 = T_25342;
  assign T_4314_74 = T_25942;
  assign T_4314_75 = T_25982;
  assign T_4314_76 = T_26202;
  assign T_4314_77 = T_25642;
  assign T_4314_78 = T_30422;
  assign T_4314_79 = T_41399;
  assign T_4314_80 = T_41527;
  assign T_4314_81 = T_41655;
  assign T_4314_82 = T_41783;
  assign T_4314_83 = T_41911;
  assign T_4314_84 = T_42039;
  assign T_4314_85 = T_42167;
  assign T_4314_86 = T_42295;
  assign T_4314_87 = T_42423;
  assign T_4314_88 = T_42551;
  assign T_4314_89 = T_42679;
  assign T_4314_90 = T_42807;
  assign T_4314_91 = T_42935;
  assign T_4314_92 = T_43063;
  assign T_4314_93 = T_43191;
  assign T_4314_94 = T_43319;
  assign T_4314_95 = T_43447;
  assign T_4314_96 = T_43575;
  assign T_4314_97 = T_43703;
  assign T_4314_98 = T_43831;
  assign T_4314_99 = T_43959;
  assign T_4314_100 = T_44087;
  assign T_4314_101 = T_44215;
  assign T_4314_102 = T_44343;
  assign T_4314_103 = T_44471;
  assign T_4314_104 = T_44599;
  assign T_4314_105 = T_44727;
  assign T_4314_106 = T_44855;
  assign T_4314_107 = T_44983;
  assign T_4314_108 = T_45111;
  assign T_4314_109 = T_45239;
  assign T_4314_110 = T_45367;
  assign T_4314_111 = T_25742;
  assign T_4314_112 = T_26182;
  assign T_4314_113 = T_25842;
  assign T_4314_114 = T_25542;
  assign T_4314_115 = T_26282;
  assign T_4314_116 = T_25442;
  assign T_4314_117 = T_26082;
  assign T_4314_118 = T_25362;
  assign T_4314_119 = T_26002;
  assign T_4314_120 = T_26262;
  assign T_4314_121 = T_45511;
  assign T_4314_122 = T_45591;
  assign T_4314_123 = T_45671;
  assign T_4314_124 = T_45751;
  assign T_4314_125 = T_45831;
  assign T_4314_126 = T_45911;
  assign T_4314_127 = T_45991;
  assign T_4314_128 = T_46071;
  assign T_4314_129 = T_46151;
  assign T_4314_130 = T_46231;
  assign T_4314_131 = T_46311;
  assign T_4314_132 = T_46391;
  assign T_4314_133 = T_46471;
  assign T_4314_134 = T_46551;
  assign T_4314_135 = T_46631;
  assign T_4314_136 = T_46711;
  assign T_4314_137 = T_46791;
  assign T_4314_138 = T_46871;
  assign T_4314_139 = T_46951;
  assign T_4314_140 = T_47031;
  assign T_4314_141 = T_25662;
  assign T_4314_142 = T_26302;
  assign T_4314_143 = T_25622;
  assign T_4314_144 = T_25922;
  assign T_4314_145 = T_25522;
  assign T_4314_146 = T_26162;
  assign T_4314_147 = T_26102;
  assign T_4314_148 = T_25822;
  assign T_4314_149 = T_25762;
  assign T_4314_150 = T_25462;
  assign T_4314_151 = T_26022;
  assign T_4314_152 = T_25902;
  assign T_4314_153 = T_26322;
  assign T_4314_154 = T_25682;
  assign T_4314_155 = T_25382;
  assign T_4314_156 = T_26242;
  assign T_4314_157 = T_25602;
  assign T_4319_0 = 1'h1;
  assign T_4319_1 = 1'h1;
  assign T_4319_2 = 1'h1;
  assign T_4319_3 = 1'h1;
  assign T_4319_4 = 1'h1;
  assign T_4319_5 = 1'h1;
  assign T_4319_6 = 1'h1;
  assign T_4319_7 = 1'h1;
  assign T_4319_8 = 1'h1;
  assign T_4319_9 = 1'h1;
  assign T_4319_10 = 1'h1;
  assign T_4319_11 = 1'h1;
  assign T_4319_12 = 1'h1;
  assign T_4319_13 = 1'h1;
  assign T_4319_14 = 1'h1;
  assign T_4319_15 = 1'h1;
  assign T_4319_16 = 1'h1;
  assign T_4319_17 = 1'h1;
  assign T_4319_18 = 1'h1;
  assign T_4319_19 = 1'h1;
  assign T_4319_20 = 1'h1;
  assign T_4319_21 = 1'h1;
  assign T_4319_22 = 1'h1;
  assign T_4319_23 = 1'h1;
  assign T_4319_24 = 1'h1;
  assign T_4319_25 = 1'h1;
  assign T_4319_26 = 1'h1;
  assign T_4319_27 = 1'h1;
  assign T_4319_28 = 1'h1;
  assign T_4319_29 = 1'h1;
  assign T_4319_30 = 1'h1;
  assign T_4319_31 = 1'h1;
  assign T_4319_32 = 1'h1;
  assign T_4319_33 = 1'h1;
  assign T_4319_34 = 1'h1;
  assign T_4319_35 = 1'h1;
  assign T_4319_36 = 1'h1;
  assign T_4319_37 = 1'h1;
  assign T_4319_38 = 1'h1;
  assign T_4319_39 = 1'h1;
  assign T_4319_40 = 1'h1;
  assign T_4319_41 = 1'h1;
  assign T_4319_42 = 1'h1;
  assign T_4319_43 = 1'h1;
  assign T_4319_44 = 1'h1;
  assign T_4319_45 = 1'h1;
  assign T_4319_46 = 1'h1;
  assign T_4319_47 = 1'h1;
  assign T_4319_48 = 1'h1;
  assign T_4319_49 = 1'h1;
  assign T_4319_50 = 1'h1;
  assign T_4319_51 = 1'h1;
  assign T_4319_52 = 1'h1;
  assign T_4319_53 = 1'h1;
  assign T_4319_54 = 1'h1;
  assign T_4319_55 = 1'h1;
  assign T_4319_56 = 1'h1;
  assign T_4319_57 = 1'h1;
  assign T_4319_58 = 1'h1;
  assign T_4319_59 = 1'h1;
  assign T_4319_60 = 1'h1;
  assign T_4319_61 = 1'h1;
  assign T_4319_62 = 1'h1;
  assign T_4319_63 = 1'h1;
  assign T_4319_64 = 1'h1;
  assign T_4319_65 = 1'h1;
  assign T_4319_66 = 1'h1;
  assign T_4319_67 = 1'h1;
  assign T_4319_68 = 1'h1;
  assign T_4319_69 = 1'h1;
  assign T_4319_70 = 1'h1;
  assign T_4319_71 = 1'h1;
  assign T_4319_72 = 1'h1;
  assign T_4319_73 = 1'h1;
  assign T_4319_74 = 1'h1;
  assign T_4319_75 = 1'h1;
  assign T_4319_76 = 1'h1;
  assign T_4319_77 = 1'h1;
  assign T_4319_78 = 1'h1;
  assign T_4319_79 = 1'h1;
  assign T_4319_80 = 1'h1;
  assign T_4319_81 = 1'h1;
  assign T_4319_82 = 1'h1;
  assign T_4319_83 = 1'h1;
  assign T_4319_84 = 1'h1;
  assign T_4319_85 = 1'h1;
  assign T_4319_86 = 1'h1;
  assign T_4319_87 = 1'h1;
  assign T_4319_88 = 1'h1;
  assign T_4319_89 = 1'h1;
  assign T_4319_90 = 1'h1;
  assign T_4319_91 = 1'h1;
  assign T_4319_92 = 1'h1;
  assign T_4319_93 = 1'h1;
  assign T_4319_94 = 1'h1;
  assign T_4319_95 = 1'h1;
  assign T_4319_96 = 1'h1;
  assign T_4319_97 = 1'h1;
  assign T_4319_98 = 1'h1;
  assign T_4319_99 = 1'h1;
  assign T_4319_100 = 1'h1;
  assign T_4319_101 = 1'h1;
  assign T_4319_102 = 1'h1;
  assign T_4319_103 = 1'h1;
  assign T_4319_104 = 1'h1;
  assign T_4319_105 = 1'h1;
  assign T_4319_106 = 1'h1;
  assign T_4319_107 = 1'h1;
  assign T_4319_108 = 1'h1;
  assign T_4319_109 = 1'h1;
  assign T_4319_110 = 1'h1;
  assign T_4319_111 = 1'h1;
  assign T_4319_112 = 1'h1;
  assign T_4319_113 = 1'h1;
  assign T_4319_114 = 1'h1;
  assign T_4319_115 = 1'h1;
  assign T_4319_116 = 1'h1;
  assign T_4319_117 = 1'h1;
  assign T_4319_118 = 1'h1;
  assign T_4319_119 = 1'h1;
  assign T_4319_120 = 1'h1;
  assign T_4319_121 = 1'h1;
  assign T_4319_122 = 1'h1;
  assign T_4319_123 = 1'h1;
  assign T_4319_124 = 1'h1;
  assign T_4319_125 = 1'h1;
  assign T_4319_126 = 1'h1;
  assign T_4319_127 = 1'h1;
  assign T_4319_128 = 1'h1;
  assign T_4319_129 = 1'h1;
  assign T_4319_130 = 1'h1;
  assign T_4319_131 = 1'h1;
  assign T_4319_132 = 1'h1;
  assign T_4319_133 = 1'h1;
  assign T_4319_134 = 1'h1;
  assign T_4319_135 = 1'h1;
  assign T_4319_136 = 1'h1;
  assign T_4319_137 = 1'h1;
  assign T_4319_138 = 1'h1;
  assign T_4319_139 = 1'h1;
  assign T_4319_140 = 1'h1;
  assign T_4319_141 = 1'h1;
  assign T_4319_142 = 1'h1;
  assign T_4319_143 = 1'h1;
  assign T_4319_144 = 1'h1;
  assign T_4319_145 = 1'h1;
  assign T_4319_146 = 1'h1;
  assign T_4319_147 = 1'h1;
  assign T_4319_148 = 1'h1;
  assign T_4319_149 = 1'h1;
  assign T_4319_150 = 1'h1;
  assign T_4319_151 = 1'h1;
  assign T_4319_152 = 1'h1;
  assign T_4319_153 = 1'h1;
  assign T_4319_154 = 1'h1;
  assign T_4319_155 = 1'h1;
  assign T_4319_156 = 1'h1;
  assign T_4319_157 = 1'h1;
  assign T_4324_0 = 1'h1;
  assign T_4324_1 = 1'h1;
  assign T_4324_2 = 1'h1;
  assign T_4324_3 = 1'h1;
  assign T_4324_4 = 1'h1;
  assign T_4324_5 = 1'h1;
  assign T_4324_6 = 1'h1;
  assign T_4324_7 = 1'h1;
  assign T_4324_8 = 1'h1;
  assign T_4324_9 = 1'h1;
  assign T_4324_10 = 1'h1;
  assign T_4324_11 = 1'h1;
  assign T_4324_12 = 1'h1;
  assign T_4324_13 = 1'h1;
  assign T_4324_14 = 1'h1;
  assign T_4324_15 = 1'h1;
  assign T_4324_16 = 1'h1;
  assign T_4324_17 = 1'h1;
  assign T_4324_18 = 1'h1;
  assign T_4324_19 = 1'h1;
  assign T_4324_20 = 1'h1;
  assign T_4324_21 = 1'h1;
  assign T_4324_22 = 1'h1;
  assign T_4324_23 = 1'h1;
  assign T_4324_24 = 1'h1;
  assign T_4324_25 = 1'h1;
  assign T_4324_26 = 1'h1;
  assign T_4324_27 = 1'h1;
  assign T_4324_28 = 1'h1;
  assign T_4324_29 = 1'h1;
  assign T_4324_30 = 1'h1;
  assign T_4324_31 = 1'h1;
  assign T_4324_32 = 1'h1;
  assign T_4324_33 = 1'h1;
  assign T_4324_34 = 1'h1;
  assign T_4324_35 = 1'h1;
  assign T_4324_36 = 1'h1;
  assign T_4324_37 = 1'h1;
  assign T_4324_38 = 1'h1;
  assign T_4324_39 = 1'h1;
  assign T_4324_40 = 1'h1;
  assign T_4324_41 = 1'h1;
  assign T_4324_42 = 1'h1;
  assign T_4324_43 = 1'h1;
  assign T_4324_44 = 1'h1;
  assign T_4324_45 = 1'h1;
  assign T_4324_46 = 1'h1;
  assign T_4324_47 = 1'h1;
  assign T_4324_48 = 1'h1;
  assign T_4324_49 = 1'h1;
  assign T_4324_50 = 1'h1;
  assign T_4324_51 = 1'h1;
  assign T_4324_52 = 1'h1;
  assign T_4324_53 = 1'h1;
  assign T_4324_54 = 1'h1;
  assign T_4324_55 = 1'h1;
  assign T_4324_56 = 1'h1;
  assign T_4324_57 = 1'h1;
  assign T_4324_58 = 1'h1;
  assign T_4324_59 = 1'h1;
  assign T_4324_60 = 1'h1;
  assign T_4324_61 = 1'h1;
  assign T_4324_62 = 1'h1;
  assign T_4324_63 = 1'h1;
  assign T_4324_64 = 1'h1;
  assign T_4324_65 = 1'h1;
  assign T_4324_66 = 1'h1;
  assign T_4324_67 = 1'h1;
  assign T_4324_68 = 1'h1;
  assign T_4324_69 = 1'h1;
  assign T_4324_70 = 1'h1;
  assign T_4324_71 = 1'h1;
  assign T_4324_72 = 1'h1;
  assign T_4324_73 = 1'h1;
  assign T_4324_74 = 1'h1;
  assign T_4324_75 = 1'h1;
  assign T_4324_76 = 1'h1;
  assign T_4324_77 = 1'h1;
  assign T_4324_78 = 1'h1;
  assign T_4324_79 = 1'h1;
  assign T_4324_80 = 1'h1;
  assign T_4324_81 = 1'h1;
  assign T_4324_82 = 1'h1;
  assign T_4324_83 = 1'h1;
  assign T_4324_84 = 1'h1;
  assign T_4324_85 = 1'h1;
  assign T_4324_86 = 1'h1;
  assign T_4324_87 = 1'h1;
  assign T_4324_88 = 1'h1;
  assign T_4324_89 = 1'h1;
  assign T_4324_90 = 1'h1;
  assign T_4324_91 = 1'h1;
  assign T_4324_92 = 1'h1;
  assign T_4324_93 = 1'h1;
  assign T_4324_94 = 1'h1;
  assign T_4324_95 = 1'h1;
  assign T_4324_96 = 1'h1;
  assign T_4324_97 = 1'h1;
  assign T_4324_98 = 1'h1;
  assign T_4324_99 = 1'h1;
  assign T_4324_100 = 1'h1;
  assign T_4324_101 = 1'h1;
  assign T_4324_102 = 1'h1;
  assign T_4324_103 = 1'h1;
  assign T_4324_104 = 1'h1;
  assign T_4324_105 = 1'h1;
  assign T_4324_106 = 1'h1;
  assign T_4324_107 = 1'h1;
  assign T_4324_108 = 1'h1;
  assign T_4324_109 = 1'h1;
  assign T_4324_110 = 1'h1;
  assign T_4324_111 = 1'h1;
  assign T_4324_112 = 1'h1;
  assign T_4324_113 = 1'h1;
  assign T_4324_114 = 1'h1;
  assign T_4324_115 = 1'h1;
  assign T_4324_116 = 1'h1;
  assign T_4324_117 = 1'h1;
  assign T_4324_118 = 1'h1;
  assign T_4324_119 = 1'h1;
  assign T_4324_120 = 1'h1;
  assign T_4324_121 = 1'h1;
  assign T_4324_122 = 1'h1;
  assign T_4324_123 = 1'h1;
  assign T_4324_124 = 1'h1;
  assign T_4324_125 = 1'h1;
  assign T_4324_126 = 1'h1;
  assign T_4324_127 = 1'h1;
  assign T_4324_128 = 1'h1;
  assign T_4324_129 = 1'h1;
  assign T_4324_130 = 1'h1;
  assign T_4324_131 = 1'h1;
  assign T_4324_132 = 1'h1;
  assign T_4324_133 = 1'h1;
  assign T_4324_134 = 1'h1;
  assign T_4324_135 = 1'h1;
  assign T_4324_136 = 1'h1;
  assign T_4324_137 = 1'h1;
  assign T_4324_138 = 1'h1;
  assign T_4324_139 = 1'h1;
  assign T_4324_140 = 1'h1;
  assign T_4324_141 = 1'h1;
  assign T_4324_142 = 1'h1;
  assign T_4324_143 = 1'h1;
  assign T_4324_144 = 1'h1;
  assign T_4324_145 = 1'h1;
  assign T_4324_146 = 1'h1;
  assign T_4324_147 = 1'h1;
  assign T_4324_148 = 1'h1;
  assign T_4324_149 = 1'h1;
  assign T_4324_150 = 1'h1;
  assign T_4324_151 = 1'h1;
  assign T_4324_152 = 1'h1;
  assign T_4324_153 = 1'h1;
  assign T_4324_154 = 1'h1;
  assign T_4324_155 = 1'h1;
  assign T_4324_156 = 1'h1;
  assign T_4324_157 = 1'h1;
  assign T_4329_0 = 1'h1;
  assign T_4329_1 = 1'h1;
  assign T_4329_2 = 1'h1;
  assign T_4329_3 = 1'h1;
  assign T_4329_4 = 1'h1;
  assign T_4329_5 = 1'h1;
  assign T_4329_6 = 1'h1;
  assign T_4329_7 = 1'h1;
  assign T_4329_8 = 1'h1;
  assign T_4329_9 = 1'h1;
  assign T_4329_10 = 1'h1;
  assign T_4329_11 = 1'h1;
  assign T_4329_12 = 1'h1;
  assign T_4329_13 = 1'h1;
  assign T_4329_14 = 1'h1;
  assign T_4329_15 = 1'h1;
  assign T_4329_16 = 1'h1;
  assign T_4329_17 = 1'h1;
  assign T_4329_18 = 1'h1;
  assign T_4329_19 = 1'h1;
  assign T_4329_20 = 1'h1;
  assign T_4329_21 = 1'h1;
  assign T_4329_22 = 1'h1;
  assign T_4329_23 = 1'h1;
  assign T_4329_24 = 1'h1;
  assign T_4329_25 = 1'h1;
  assign T_4329_26 = 1'h1;
  assign T_4329_27 = 1'h1;
  assign T_4329_28 = 1'h1;
  assign T_4329_29 = 1'h1;
  assign T_4329_30 = 1'h1;
  assign T_4329_31 = 1'h1;
  assign T_4329_32 = 1'h1;
  assign T_4329_33 = 1'h1;
  assign T_4329_34 = 1'h1;
  assign T_4329_35 = 1'h1;
  assign T_4329_36 = 1'h1;
  assign T_4329_37 = 1'h1;
  assign T_4329_38 = 1'h1;
  assign T_4329_39 = 1'h1;
  assign T_4329_40 = 1'h1;
  assign T_4329_41 = 1'h1;
  assign T_4329_42 = 1'h1;
  assign T_4329_43 = 1'h1;
  assign T_4329_44 = 1'h1;
  assign T_4329_45 = 1'h1;
  assign T_4329_46 = 1'h1;
  assign T_4329_47 = 1'h1;
  assign T_4329_48 = 1'h1;
  assign T_4329_49 = 1'h1;
  assign T_4329_50 = 1'h1;
  assign T_4329_51 = 1'h1;
  assign T_4329_52 = 1'h1;
  assign T_4329_53 = 1'h1;
  assign T_4329_54 = 1'h1;
  assign T_4329_55 = 1'h1;
  assign T_4329_56 = 1'h1;
  assign T_4329_57 = 1'h1;
  assign T_4329_58 = 1'h1;
  assign T_4329_59 = 1'h1;
  assign T_4329_60 = 1'h1;
  assign T_4329_61 = 1'h1;
  assign T_4329_62 = 1'h1;
  assign T_4329_63 = 1'h1;
  assign T_4329_64 = 1'h1;
  assign T_4329_65 = 1'h1;
  assign T_4329_66 = 1'h1;
  assign T_4329_67 = 1'h1;
  assign T_4329_68 = 1'h1;
  assign T_4329_69 = 1'h1;
  assign T_4329_70 = 1'h1;
  assign T_4329_71 = 1'h1;
  assign T_4329_72 = 1'h1;
  assign T_4329_73 = 1'h1;
  assign T_4329_74 = 1'h1;
  assign T_4329_75 = 1'h1;
  assign T_4329_76 = 1'h1;
  assign T_4329_77 = 1'h1;
  assign T_4329_78 = 1'h1;
  assign T_4329_79 = 1'h1;
  assign T_4329_80 = 1'h1;
  assign T_4329_81 = 1'h1;
  assign T_4329_82 = 1'h1;
  assign T_4329_83 = 1'h1;
  assign T_4329_84 = 1'h1;
  assign T_4329_85 = 1'h1;
  assign T_4329_86 = 1'h1;
  assign T_4329_87 = 1'h1;
  assign T_4329_88 = 1'h1;
  assign T_4329_89 = 1'h1;
  assign T_4329_90 = 1'h1;
  assign T_4329_91 = 1'h1;
  assign T_4329_92 = 1'h1;
  assign T_4329_93 = 1'h1;
  assign T_4329_94 = 1'h1;
  assign T_4329_95 = 1'h1;
  assign T_4329_96 = 1'h1;
  assign T_4329_97 = 1'h1;
  assign T_4329_98 = 1'h1;
  assign T_4329_99 = 1'h1;
  assign T_4329_100 = 1'h1;
  assign T_4329_101 = 1'h1;
  assign T_4329_102 = 1'h1;
  assign T_4329_103 = 1'h1;
  assign T_4329_104 = 1'h1;
  assign T_4329_105 = 1'h1;
  assign T_4329_106 = 1'h1;
  assign T_4329_107 = 1'h1;
  assign T_4329_108 = 1'h1;
  assign T_4329_109 = 1'h1;
  assign T_4329_110 = 1'h1;
  assign T_4329_111 = 1'h1;
  assign T_4329_112 = 1'h1;
  assign T_4329_113 = 1'h1;
  assign T_4329_114 = 1'h1;
  assign T_4329_115 = 1'h1;
  assign T_4329_116 = 1'h1;
  assign T_4329_117 = 1'h1;
  assign T_4329_118 = 1'h1;
  assign T_4329_119 = 1'h1;
  assign T_4329_120 = 1'h1;
  assign T_4329_121 = 1'h1;
  assign T_4329_122 = 1'h1;
  assign T_4329_123 = 1'h1;
  assign T_4329_124 = 1'h1;
  assign T_4329_125 = 1'h1;
  assign T_4329_126 = 1'h1;
  assign T_4329_127 = 1'h1;
  assign T_4329_128 = 1'h1;
  assign T_4329_129 = 1'h1;
  assign T_4329_130 = 1'h1;
  assign T_4329_131 = 1'h1;
  assign T_4329_132 = 1'h1;
  assign T_4329_133 = 1'h1;
  assign T_4329_134 = 1'h1;
  assign T_4329_135 = 1'h1;
  assign T_4329_136 = 1'h1;
  assign T_4329_137 = 1'h1;
  assign T_4329_138 = 1'h1;
  assign T_4329_139 = 1'h1;
  assign T_4329_140 = 1'h1;
  assign T_4329_141 = 1'h1;
  assign T_4329_142 = 1'h1;
  assign T_4329_143 = 1'h1;
  assign T_4329_144 = 1'h1;
  assign T_4329_145 = 1'h1;
  assign T_4329_146 = 1'h1;
  assign T_4329_147 = 1'h1;
  assign T_4329_148 = 1'h1;
  assign T_4329_149 = 1'h1;
  assign T_4329_150 = 1'h1;
  assign T_4329_151 = 1'h1;
  assign T_4329_152 = 1'h1;
  assign T_4329_153 = 1'h1;
  assign T_4329_154 = 1'h1;
  assign T_4329_155 = 1'h1;
  assign T_4329_156 = 1'h1;
  assign T_4329_157 = 1'h1;
  assign T_4334_0 = 1'h1;
  assign T_4334_1 = 1'h1;
  assign T_4334_2 = 1'h1;
  assign T_4334_3 = 1'h1;
  assign T_4334_4 = 1'h1;
  assign T_4334_5 = 1'h1;
  assign T_4334_6 = 1'h1;
  assign T_4334_7 = 1'h1;
  assign T_4334_8 = 1'h1;
  assign T_4334_9 = 1'h1;
  assign T_4334_10 = 1'h1;
  assign T_4334_11 = 1'h1;
  assign T_4334_12 = 1'h1;
  assign T_4334_13 = 1'h1;
  assign T_4334_14 = 1'h1;
  assign T_4334_15 = 1'h1;
  assign T_4334_16 = 1'h1;
  assign T_4334_17 = 1'h1;
  assign T_4334_18 = 1'h1;
  assign T_4334_19 = 1'h1;
  assign T_4334_20 = 1'h1;
  assign T_4334_21 = 1'h1;
  assign T_4334_22 = 1'h1;
  assign T_4334_23 = 1'h1;
  assign T_4334_24 = 1'h1;
  assign T_4334_25 = 1'h1;
  assign T_4334_26 = 1'h1;
  assign T_4334_27 = 1'h1;
  assign T_4334_28 = 1'h1;
  assign T_4334_29 = 1'h1;
  assign T_4334_30 = 1'h1;
  assign T_4334_31 = 1'h1;
  assign T_4334_32 = 1'h1;
  assign T_4334_33 = 1'h1;
  assign T_4334_34 = 1'h1;
  assign T_4334_35 = 1'h1;
  assign T_4334_36 = 1'h1;
  assign T_4334_37 = 1'h1;
  assign T_4334_38 = 1'h1;
  assign T_4334_39 = 1'h1;
  assign T_4334_40 = 1'h1;
  assign T_4334_41 = 1'h1;
  assign T_4334_42 = 1'h1;
  assign T_4334_43 = 1'h1;
  assign T_4334_44 = 1'h1;
  assign T_4334_45 = 1'h1;
  assign T_4334_46 = 1'h1;
  assign T_4334_47 = 1'h1;
  assign T_4334_48 = 1'h1;
  assign T_4334_49 = 1'h1;
  assign T_4334_50 = 1'h1;
  assign T_4334_51 = 1'h1;
  assign T_4334_52 = 1'h1;
  assign T_4334_53 = 1'h1;
  assign T_4334_54 = 1'h1;
  assign T_4334_55 = 1'h1;
  assign T_4334_56 = 1'h1;
  assign T_4334_57 = 1'h1;
  assign T_4334_58 = 1'h1;
  assign T_4334_59 = 1'h1;
  assign T_4334_60 = 1'h1;
  assign T_4334_61 = 1'h1;
  assign T_4334_62 = 1'h1;
  assign T_4334_63 = 1'h1;
  assign T_4334_64 = 1'h1;
  assign T_4334_65 = 1'h1;
  assign T_4334_66 = 1'h1;
  assign T_4334_67 = 1'h1;
  assign T_4334_68 = 1'h1;
  assign T_4334_69 = 1'h1;
  assign T_4334_70 = 1'h1;
  assign T_4334_71 = 1'h1;
  assign T_4334_72 = 1'h1;
  assign T_4334_73 = 1'h1;
  assign T_4334_74 = 1'h1;
  assign T_4334_75 = 1'h1;
  assign T_4334_76 = 1'h1;
  assign T_4334_77 = 1'h1;
  assign T_4334_78 = 1'h1;
  assign T_4334_79 = 1'h1;
  assign T_4334_80 = 1'h1;
  assign T_4334_81 = 1'h1;
  assign T_4334_82 = 1'h1;
  assign T_4334_83 = 1'h1;
  assign T_4334_84 = 1'h1;
  assign T_4334_85 = 1'h1;
  assign T_4334_86 = 1'h1;
  assign T_4334_87 = 1'h1;
  assign T_4334_88 = 1'h1;
  assign T_4334_89 = 1'h1;
  assign T_4334_90 = 1'h1;
  assign T_4334_91 = 1'h1;
  assign T_4334_92 = 1'h1;
  assign T_4334_93 = 1'h1;
  assign T_4334_94 = 1'h1;
  assign T_4334_95 = 1'h1;
  assign T_4334_96 = 1'h1;
  assign T_4334_97 = 1'h1;
  assign T_4334_98 = 1'h1;
  assign T_4334_99 = 1'h1;
  assign T_4334_100 = 1'h1;
  assign T_4334_101 = 1'h1;
  assign T_4334_102 = 1'h1;
  assign T_4334_103 = 1'h1;
  assign T_4334_104 = 1'h1;
  assign T_4334_105 = 1'h1;
  assign T_4334_106 = 1'h1;
  assign T_4334_107 = 1'h1;
  assign T_4334_108 = 1'h1;
  assign T_4334_109 = 1'h1;
  assign T_4334_110 = 1'h1;
  assign T_4334_111 = 1'h1;
  assign T_4334_112 = 1'h1;
  assign T_4334_113 = 1'h1;
  assign T_4334_114 = 1'h1;
  assign T_4334_115 = 1'h1;
  assign T_4334_116 = 1'h1;
  assign T_4334_117 = 1'h1;
  assign T_4334_118 = 1'h1;
  assign T_4334_119 = 1'h1;
  assign T_4334_120 = 1'h1;
  assign T_4334_121 = 1'h1;
  assign T_4334_122 = 1'h1;
  assign T_4334_123 = 1'h1;
  assign T_4334_124 = 1'h1;
  assign T_4334_125 = 1'h1;
  assign T_4334_126 = 1'h1;
  assign T_4334_127 = 1'h1;
  assign T_4334_128 = 1'h1;
  assign T_4334_129 = 1'h1;
  assign T_4334_130 = 1'h1;
  assign T_4334_131 = 1'h1;
  assign T_4334_132 = 1'h1;
  assign T_4334_133 = 1'h1;
  assign T_4334_134 = 1'h1;
  assign T_4334_135 = 1'h1;
  assign T_4334_136 = 1'h1;
  assign T_4334_137 = 1'h1;
  assign T_4334_138 = 1'h1;
  assign T_4334_139 = 1'h1;
  assign T_4334_140 = 1'h1;
  assign T_4334_141 = 1'h1;
  assign T_4334_142 = 1'h1;
  assign T_4334_143 = 1'h1;
  assign T_4334_144 = 1'h1;
  assign T_4334_145 = 1'h1;
  assign T_4334_146 = 1'h1;
  assign T_4334_147 = 1'h1;
  assign T_4334_148 = 1'h1;
  assign T_4334_149 = 1'h1;
  assign T_4334_150 = 1'h1;
  assign T_4334_151 = 1'h1;
  assign T_4334_152 = 1'h1;
  assign T_4334_153 = 1'h1;
  assign T_4334_154 = 1'h1;
  assign T_4334_155 = 1'h1;
  assign T_4334_156 = 1'h1;
  assign T_4334_157 = 1'h1;
  assign T_4339_0 = T_35627;
  assign T_4339_1 = T_35755;
  assign T_4339_2 = T_35883;
  assign T_4339_3 = T_36011;
  assign T_4339_4 = T_36139;
  assign T_4339_5 = T_36267;
  assign T_4339_6 = T_36395;
  assign T_4339_7 = T_36523;
  assign T_4339_8 = T_36651;
  assign T_4339_9 = T_36779;
  assign T_4339_10 = T_36907;
  assign T_4339_11 = T_37035;
  assign T_4339_12 = T_37163;
  assign T_4339_13 = T_37291;
  assign T_4339_14 = T_37419;
  assign T_4339_15 = T_37547;
  assign T_4339_16 = T_37675;
  assign T_4339_17 = T_37803;
  assign T_4339_18 = T_37931;
  assign T_4339_19 = T_38059;
  assign T_4339_20 = T_38187;
  assign T_4339_21 = T_38315;
  assign T_4339_22 = T_38443;
  assign T_4339_23 = T_38571;
  assign T_4339_24 = T_38699;
  assign T_4339_25 = T_38827;
  assign T_4339_26 = T_38955;
  assign T_4339_27 = T_39083;
  assign T_4339_28 = T_39211;
  assign T_4339_29 = T_39339;
  assign T_4339_30 = T_39467;
  assign T_4339_31 = T_39595;
  assign T_4339_32 = T_25306;
  assign T_4339_33 = T_25406;
  assign T_4339_34 = T_25506;
  assign T_4339_35 = T_26146;
  assign T_4339_36 = T_25786;
  assign T_4339_37 = T_26046;
  assign T_4339_38 = T_25806;
  assign T_4339_39 = T_25586;
  assign T_4339_40 = T_25706;
  assign T_4339_41 = T_39723;
  assign T_4339_42 = T_39803;
  assign T_4339_43 = T_39883;
  assign T_4339_44 = T_39963;
  assign T_4339_45 = T_40043;
  assign T_4339_46 = T_40123;
  assign T_4339_47 = T_40203;
  assign T_4339_48 = T_40283;
  assign T_4339_49 = T_40363;
  assign T_4339_50 = T_40443;
  assign T_4339_51 = T_40523;
  assign T_4339_52 = T_40603;
  assign T_4339_53 = T_40683;
  assign T_4339_54 = T_40763;
  assign T_4339_55 = T_40843;
  assign T_4339_56 = T_40923;
  assign T_4339_57 = T_41003;
  assign T_4339_58 = T_41083;
  assign T_4339_59 = T_41163;
  assign T_4339_60 = T_41243;
  assign T_4339_61 = T_26226;
  assign T_4339_62 = T_25886;
  assign T_4339_63 = T_30446;
  assign T_4339_64 = T_25326;
  assign T_4339_65 = T_25426;
  assign T_4339_66 = T_25866;
  assign T_4339_67 = T_26066;
  assign T_4339_68 = T_25726;
  assign T_4339_69 = T_25966;
  assign T_4339_70 = T_25486;
  assign T_4339_71 = T_25566;
  assign T_4339_72 = T_26126;
  assign T_4339_73 = T_25346;
  assign T_4339_74 = T_25946;
  assign T_4339_75 = T_25986;
  assign T_4339_76 = T_26206;
  assign T_4339_77 = T_25646;
  assign T_4339_78 = T_30426;
  assign T_4339_79 = T_41431;
  assign T_4339_80 = T_41559;
  assign T_4339_81 = T_41687;
  assign T_4339_82 = T_41815;
  assign T_4339_83 = T_41943;
  assign T_4339_84 = T_42071;
  assign T_4339_85 = T_42199;
  assign T_4339_86 = T_42327;
  assign T_4339_87 = T_42455;
  assign T_4339_88 = T_42583;
  assign T_4339_89 = T_42711;
  assign T_4339_90 = T_42839;
  assign T_4339_91 = T_42967;
  assign T_4339_92 = T_43095;
  assign T_4339_93 = T_43223;
  assign T_4339_94 = T_43351;
  assign T_4339_95 = T_43479;
  assign T_4339_96 = T_43607;
  assign T_4339_97 = T_43735;
  assign T_4339_98 = T_43863;
  assign T_4339_99 = T_43991;
  assign T_4339_100 = T_44119;
  assign T_4339_101 = T_44247;
  assign T_4339_102 = T_44375;
  assign T_4339_103 = T_44503;
  assign T_4339_104 = T_44631;
  assign T_4339_105 = T_44759;
  assign T_4339_106 = T_44887;
  assign T_4339_107 = T_45015;
  assign T_4339_108 = T_45143;
  assign T_4339_109 = T_45271;
  assign T_4339_110 = T_45399;
  assign T_4339_111 = T_25746;
  assign T_4339_112 = T_26186;
  assign T_4339_113 = T_25846;
  assign T_4339_114 = T_25546;
  assign T_4339_115 = T_26286;
  assign T_4339_116 = T_25446;
  assign T_4339_117 = T_26086;
  assign T_4339_118 = T_25366;
  assign T_4339_119 = T_26006;
  assign T_4339_120 = T_26266;
  assign T_4339_121 = T_45531;
  assign T_4339_122 = T_45611;
  assign T_4339_123 = T_45691;
  assign T_4339_124 = T_45771;
  assign T_4339_125 = T_45851;
  assign T_4339_126 = T_45931;
  assign T_4339_127 = T_46011;
  assign T_4339_128 = T_46091;
  assign T_4339_129 = T_46171;
  assign T_4339_130 = T_46251;
  assign T_4339_131 = T_46331;
  assign T_4339_132 = T_46411;
  assign T_4339_133 = T_46491;
  assign T_4339_134 = T_46571;
  assign T_4339_135 = T_46651;
  assign T_4339_136 = T_46731;
  assign T_4339_137 = T_46811;
  assign T_4339_138 = T_46891;
  assign T_4339_139 = T_46971;
  assign T_4339_140 = T_47051;
  assign T_4339_141 = T_25666;
  assign T_4339_142 = T_26306;
  assign T_4339_143 = T_25626;
  assign T_4339_144 = T_25926;
  assign T_4339_145 = T_25526;
  assign T_4339_146 = T_26166;
  assign T_4339_147 = T_26106;
  assign T_4339_148 = T_25826;
  assign T_4339_149 = T_25766;
  assign T_4339_150 = T_25466;
  assign T_4339_151 = T_26026;
  assign T_4339_152 = T_25906;
  assign T_4339_153 = T_26326;
  assign T_4339_154 = T_25686;
  assign T_4339_155 = T_25386;
  assign T_4339_156 = T_26246;
  assign T_4339_157 = T_25606;
  assign T_4344_0 = T_35659;
  assign T_4344_1 = T_35787;
  assign T_4344_2 = T_35915;
  assign T_4344_3 = T_36043;
  assign T_4344_4 = T_36171;
  assign T_4344_5 = T_36299;
  assign T_4344_6 = T_36427;
  assign T_4344_7 = T_36555;
  assign T_4344_8 = T_36683;
  assign T_4344_9 = T_36811;
  assign T_4344_10 = T_36939;
  assign T_4344_11 = T_37067;
  assign T_4344_12 = T_37195;
  assign T_4344_13 = T_37323;
  assign T_4344_14 = T_37451;
  assign T_4344_15 = T_37579;
  assign T_4344_16 = T_37707;
  assign T_4344_17 = T_37835;
  assign T_4344_18 = T_37963;
  assign T_4344_19 = T_38091;
  assign T_4344_20 = T_38219;
  assign T_4344_21 = T_38347;
  assign T_4344_22 = T_38475;
  assign T_4344_23 = T_38603;
  assign T_4344_24 = T_38731;
  assign T_4344_25 = T_38859;
  assign T_4344_26 = T_38987;
  assign T_4344_27 = T_39115;
  assign T_4344_28 = T_39243;
  assign T_4344_29 = T_39371;
  assign T_4344_30 = T_39499;
  assign T_4344_31 = T_39627;
  assign T_4344_32 = T_25312;
  assign T_4344_33 = T_25412;
  assign T_4344_34 = T_25512;
  assign T_4344_35 = T_26152;
  assign T_4344_36 = T_25792;
  assign T_4344_37 = T_26052;
  assign T_4344_38 = T_25812;
  assign T_4344_39 = T_25592;
  assign T_4344_40 = T_25712;
  assign T_4344_41 = T_39743;
  assign T_4344_42 = T_39823;
  assign T_4344_43 = T_39903;
  assign T_4344_44 = T_39983;
  assign T_4344_45 = T_40063;
  assign T_4344_46 = T_40143;
  assign T_4344_47 = T_40223;
  assign T_4344_48 = T_40303;
  assign T_4344_49 = T_40383;
  assign T_4344_50 = T_40463;
  assign T_4344_51 = T_40543;
  assign T_4344_52 = T_40623;
  assign T_4344_53 = T_40703;
  assign T_4344_54 = T_40783;
  assign T_4344_55 = T_40863;
  assign T_4344_56 = T_40943;
  assign T_4344_57 = T_41023;
  assign T_4344_58 = T_41103;
  assign T_4344_59 = T_41183;
  assign T_4344_60 = T_41263;
  assign T_4344_61 = T_26232;
  assign T_4344_62 = T_25892;
  assign T_4344_63 = T_30452;
  assign T_4344_64 = T_25332;
  assign T_4344_65 = T_25432;
  assign T_4344_66 = T_25872;
  assign T_4344_67 = T_26072;
  assign T_4344_68 = T_25732;
  assign T_4344_69 = T_25972;
  assign T_4344_70 = T_25492;
  assign T_4344_71 = T_25572;
  assign T_4344_72 = T_26132;
  assign T_4344_73 = T_25352;
  assign T_4344_74 = T_25952;
  assign T_4344_75 = T_25992;
  assign T_4344_76 = T_26212;
  assign T_4344_77 = T_25652;
  assign T_4344_78 = T_30432;
  assign T_4344_79 = T_41463;
  assign T_4344_80 = T_41591;
  assign T_4344_81 = T_41719;
  assign T_4344_82 = T_41847;
  assign T_4344_83 = T_41975;
  assign T_4344_84 = T_42103;
  assign T_4344_85 = T_42231;
  assign T_4344_86 = T_42359;
  assign T_4344_87 = T_42487;
  assign T_4344_88 = T_42615;
  assign T_4344_89 = T_42743;
  assign T_4344_90 = T_42871;
  assign T_4344_91 = T_42999;
  assign T_4344_92 = T_43127;
  assign T_4344_93 = T_43255;
  assign T_4344_94 = T_43383;
  assign T_4344_95 = T_43511;
  assign T_4344_96 = T_43639;
  assign T_4344_97 = T_43767;
  assign T_4344_98 = T_43895;
  assign T_4344_99 = T_44023;
  assign T_4344_100 = T_44151;
  assign T_4344_101 = T_44279;
  assign T_4344_102 = T_44407;
  assign T_4344_103 = T_44535;
  assign T_4344_104 = T_44663;
  assign T_4344_105 = T_44791;
  assign T_4344_106 = T_44919;
  assign T_4344_107 = T_45047;
  assign T_4344_108 = T_45175;
  assign T_4344_109 = T_45303;
  assign T_4344_110 = T_45431;
  assign T_4344_111 = T_25752;
  assign T_4344_112 = T_26192;
  assign T_4344_113 = T_25852;
  assign T_4344_114 = T_25552;
  assign T_4344_115 = T_26292;
  assign T_4344_116 = T_25452;
  assign T_4344_117 = T_26092;
  assign T_4344_118 = T_25372;
  assign T_4344_119 = T_26012;
  assign T_4344_120 = T_26272;
  assign T_4344_121 = T_45551;
  assign T_4344_122 = T_45631;
  assign T_4344_123 = T_45711;
  assign T_4344_124 = T_45791;
  assign T_4344_125 = T_45871;
  assign T_4344_126 = T_45951;
  assign T_4344_127 = T_46031;
  assign T_4344_128 = T_46111;
  assign T_4344_129 = T_46191;
  assign T_4344_130 = T_46271;
  assign T_4344_131 = T_46351;
  assign T_4344_132 = T_46431;
  assign T_4344_133 = T_46511;
  assign T_4344_134 = T_46591;
  assign T_4344_135 = T_46671;
  assign T_4344_136 = T_46751;
  assign T_4344_137 = T_46831;
  assign T_4344_138 = T_46911;
  assign T_4344_139 = T_46991;
  assign T_4344_140 = T_47071;
  assign T_4344_141 = T_25672;
  assign T_4344_142 = T_26312;
  assign T_4344_143 = T_25632;
  assign T_4344_144 = T_25932;
  assign T_4344_145 = T_25532;
  assign T_4344_146 = T_26172;
  assign T_4344_147 = T_26112;
  assign T_4344_148 = T_25832;
  assign T_4344_149 = T_25772;
  assign T_4344_150 = T_25472;
  assign T_4344_151 = T_26032;
  assign T_4344_152 = T_25912;
  assign T_4344_153 = T_26332;
  assign T_4344_154 = T_25692;
  assign T_4344_155 = T_25392;
  assign T_4344_156 = T_26252;
  assign T_4344_157 = T_25612;
  assign T_6906 = T_3205_bits_mask[0];
  assign T_6907 = T_3205_bits_mask[1];
  assign T_6908 = T_3205_bits_mask[2];
  assign T_6909 = T_3205_bits_mask[3];
  assign T_6913 = T_6906 ? 8'hff : 8'h0;
  assign T_6917 = T_6907 ? 8'hff : 8'h0;
  assign T_6921 = T_6908 ? 8'hff : 8'h0;
  assign T_6925 = T_6909 ? 8'hff : 8'h0;
  assign T_6926 = {T_6917,T_6913};
  assign T_6927 = {T_6925,T_6921};
  assign T_6928 = {T_6927,T_6926};
  assign T_6952 = T_6928[0];
  assign T_6956 = ~ T_6952;
  assign T_6958 = T_6956 == 1'h0;
  assign T_6972 = T_3205_bits_data[0];
  assign T_6992 = T_6928[1];
  assign T_6996 = ~ T_6992;
  assign T_6998 = T_6996 == 1'h0;
  assign T_7012 = T_3205_bits_data[1];
  assign GEN_3514 = {{1'd0}, pending_1};
  assign T_7027 = GEN_3514 << 1;
  assign GEN_3515 = {{1'd0}, pending_0};
  assign T_7031 = GEN_3515 | T_7027;
  assign T_7032 = T_6928[2];
  assign T_7036 = ~ T_7032;
  assign T_7038 = T_7036 == 1'h0;
  assign T_7052 = T_3205_bits_data[2];
  assign GEN_3516 = {{2'd0}, pending_2};
  assign T_7067 = GEN_3516 << 2;
  assign GEN_3517 = {{1'd0}, T_7031};
  assign T_7071 = GEN_3517 | T_7067;
  assign T_7072 = T_6928[3];
  assign T_7076 = ~ T_7072;
  assign T_7078 = T_7076 == 1'h0;
  assign T_7092 = T_3205_bits_data[3];
  assign GEN_3518 = {{3'd0}, pending_3};
  assign T_7107 = GEN_3518 << 3;
  assign GEN_3519 = {{1'd0}, T_7071};
  assign T_7111 = GEN_3519 | T_7107;
  assign T_7112 = T_6928[4];
  assign T_7116 = ~ T_7112;
  assign T_7118 = T_7116 == 1'h0;
  assign T_7132 = T_3205_bits_data[4];
  assign GEN_3520 = {{4'd0}, pending_4};
  assign T_7147 = GEN_3520 << 4;
  assign GEN_3521 = {{1'd0}, T_7111};
  assign T_7151 = GEN_3521 | T_7147;
  assign T_7152 = T_6928[5];
  assign T_7156 = ~ T_7152;
  assign T_7158 = T_7156 == 1'h0;
  assign T_7172 = T_3205_bits_data[5];
  assign GEN_3522 = {{5'd0}, pending_5};
  assign T_7187 = GEN_3522 << 5;
  assign GEN_3523 = {{1'd0}, T_7151};
  assign T_7191 = GEN_3523 | T_7187;
  assign T_7192 = T_6928[6];
  assign T_7196 = ~ T_7192;
  assign T_7198 = T_7196 == 1'h0;
  assign T_7212 = T_3205_bits_data[6];
  assign GEN_3524 = {{6'd0}, pending_6};
  assign T_7227 = GEN_3524 << 6;
  assign GEN_3525 = {{1'd0}, T_7191};
  assign T_7231 = GEN_3525 | T_7227;
  assign T_7232 = T_6928[7];
  assign T_7236 = ~ T_7232;
  assign T_7238 = T_7236 == 1'h0;
  assign T_7252 = T_3205_bits_data[7];
  assign GEN_3526 = {{7'd0}, pending_7};
  assign T_7267 = GEN_3526 << 7;
  assign GEN_3527 = {{1'd0}, T_7231};
  assign T_7271 = GEN_3527 | T_7267;
  assign T_7272 = T_6928[8];
  assign T_7276 = ~ T_7272;
  assign T_7278 = T_7276 == 1'h0;
  assign T_7292 = T_3205_bits_data[8];
  assign GEN_3528 = {{8'd0}, pending_8};
  assign T_7307 = GEN_3528 << 8;
  assign GEN_3529 = {{1'd0}, T_7271};
  assign T_7311 = GEN_3529 | T_7307;
  assign T_7312 = T_6928[9];
  assign T_7316 = ~ T_7312;
  assign T_7318 = T_7316 == 1'h0;
  assign T_7332 = T_3205_bits_data[9];
  assign GEN_3530 = {{9'd0}, pending_9};
  assign T_7347 = GEN_3530 << 9;
  assign GEN_3531 = {{1'd0}, T_7311};
  assign T_7351 = GEN_3531 | T_7347;
  assign T_7352 = T_6928[10];
  assign T_7356 = ~ T_7352;
  assign T_7358 = T_7356 == 1'h0;
  assign T_7372 = T_3205_bits_data[10];
  assign GEN_3532 = {{10'd0}, pending_10};
  assign T_7387 = GEN_3532 << 10;
  assign GEN_3533 = {{1'd0}, T_7351};
  assign T_7391 = GEN_3533 | T_7387;
  assign T_7392 = T_6928[11];
  assign T_7396 = ~ T_7392;
  assign T_7398 = T_7396 == 1'h0;
  assign T_7412 = T_3205_bits_data[11];
  assign GEN_3534 = {{11'd0}, pending_11};
  assign T_7427 = GEN_3534 << 11;
  assign GEN_3535 = {{1'd0}, T_7391};
  assign T_7431 = GEN_3535 | T_7427;
  assign T_7432 = T_6928[12];
  assign T_7436 = ~ T_7432;
  assign T_7438 = T_7436 == 1'h0;
  assign T_7452 = T_3205_bits_data[12];
  assign GEN_3536 = {{12'd0}, pending_12};
  assign T_7467 = GEN_3536 << 12;
  assign GEN_3537 = {{1'd0}, T_7431};
  assign T_7471 = GEN_3537 | T_7467;
  assign T_7472 = T_6928[13];
  assign T_7476 = ~ T_7472;
  assign T_7478 = T_7476 == 1'h0;
  assign T_7492 = T_3205_bits_data[13];
  assign GEN_3538 = {{13'd0}, pending_13};
  assign T_7507 = GEN_3538 << 13;
  assign GEN_3539 = {{1'd0}, T_7471};
  assign T_7511 = GEN_3539 | T_7507;
  assign T_7512 = T_6928[14];
  assign T_7516 = ~ T_7512;
  assign T_7518 = T_7516 == 1'h0;
  assign T_7532 = T_3205_bits_data[14];
  assign GEN_3540 = {{14'd0}, pending_14};
  assign T_7547 = GEN_3540 << 14;
  assign GEN_3541 = {{1'd0}, T_7511};
  assign T_7551 = GEN_3541 | T_7547;
  assign T_7552 = T_6928[15];
  assign T_7556 = ~ T_7552;
  assign T_7558 = T_7556 == 1'h0;
  assign T_7572 = T_3205_bits_data[15];
  assign GEN_3542 = {{15'd0}, pending_15};
  assign T_7587 = GEN_3542 << 15;
  assign GEN_3543 = {{1'd0}, T_7551};
  assign T_7591 = GEN_3543 | T_7587;
  assign T_7592 = T_6928[16];
  assign T_7596 = ~ T_7592;
  assign T_7598 = T_7596 == 1'h0;
  assign T_7612 = T_3205_bits_data[16];
  assign GEN_3544 = {{16'd0}, pending_16};
  assign T_7627 = GEN_3544 << 16;
  assign GEN_3545 = {{1'd0}, T_7591};
  assign T_7631 = GEN_3545 | T_7627;
  assign T_7632 = T_6928[17];
  assign T_7636 = ~ T_7632;
  assign T_7638 = T_7636 == 1'h0;
  assign T_7652 = T_3205_bits_data[17];
  assign GEN_3546 = {{17'd0}, pending_17};
  assign T_7667 = GEN_3546 << 17;
  assign GEN_3547 = {{1'd0}, T_7631};
  assign T_7671 = GEN_3547 | T_7667;
  assign T_7672 = T_6928[18];
  assign T_7676 = ~ T_7672;
  assign T_7678 = T_7676 == 1'h0;
  assign T_7692 = T_3205_bits_data[18];
  assign GEN_3548 = {{18'd0}, pending_18};
  assign T_7707 = GEN_3548 << 18;
  assign GEN_3549 = {{1'd0}, T_7671};
  assign T_7711 = GEN_3549 | T_7707;
  assign T_7712 = T_6928[19];
  assign T_7716 = ~ T_7712;
  assign T_7718 = T_7716 == 1'h0;
  assign T_7732 = T_3205_bits_data[19];
  assign GEN_3550 = {{19'd0}, pending_19};
  assign T_7747 = GEN_3550 << 19;
  assign GEN_3551 = {{1'd0}, T_7711};
  assign T_7751 = GEN_3551 | T_7747;
  assign T_7752 = T_6928[20];
  assign T_7756 = ~ T_7752;
  assign T_7758 = T_7756 == 1'h0;
  assign T_7772 = T_3205_bits_data[20];
  assign GEN_3552 = {{20'd0}, pending_20};
  assign T_7787 = GEN_3552 << 20;
  assign GEN_3553 = {{1'd0}, T_7751};
  assign T_7791 = GEN_3553 | T_7787;
  assign T_7792 = T_6928[21];
  assign T_7796 = ~ T_7792;
  assign T_7798 = T_7796 == 1'h0;
  assign T_7812 = T_3205_bits_data[21];
  assign GEN_3554 = {{21'd0}, pending_21};
  assign T_7827 = GEN_3554 << 21;
  assign GEN_3555 = {{1'd0}, T_7791};
  assign T_7831 = GEN_3555 | T_7827;
  assign T_7832 = T_6928[22];
  assign T_7836 = ~ T_7832;
  assign T_7838 = T_7836 == 1'h0;
  assign T_7852 = T_3205_bits_data[22];
  assign GEN_3556 = {{22'd0}, pending_22};
  assign T_7867 = GEN_3556 << 22;
  assign GEN_3557 = {{1'd0}, T_7831};
  assign T_7871 = GEN_3557 | T_7867;
  assign T_7872 = T_6928[23];
  assign T_7876 = ~ T_7872;
  assign T_7878 = T_7876 == 1'h0;
  assign T_7892 = T_3205_bits_data[23];
  assign GEN_3558 = {{23'd0}, pending_23};
  assign T_7907 = GEN_3558 << 23;
  assign GEN_3559 = {{1'd0}, T_7871};
  assign T_7911 = GEN_3559 | T_7907;
  assign T_7912 = T_6928[24];
  assign T_7916 = ~ T_7912;
  assign T_7918 = T_7916 == 1'h0;
  assign T_7932 = T_3205_bits_data[24];
  assign GEN_3560 = {{24'd0}, pending_24};
  assign T_7947 = GEN_3560 << 24;
  assign GEN_3561 = {{1'd0}, T_7911};
  assign T_7951 = GEN_3561 | T_7947;
  assign T_7952 = T_6928[25];
  assign T_7956 = ~ T_7952;
  assign T_7958 = T_7956 == 1'h0;
  assign T_7972 = T_3205_bits_data[25];
  assign GEN_3562 = {{25'd0}, pending_25};
  assign T_7987 = GEN_3562 << 25;
  assign GEN_3563 = {{1'd0}, T_7951};
  assign T_7991 = GEN_3563 | T_7987;
  assign T_7992 = T_6928[26];
  assign T_7996 = ~ T_7992;
  assign T_7998 = T_7996 == 1'h0;
  assign T_8012 = T_3205_bits_data[26];
  assign GEN_3564 = {{26'd0}, pending_26};
  assign T_8027 = GEN_3564 << 26;
  assign GEN_3565 = {{1'd0}, T_7991};
  assign T_8031 = GEN_3565 | T_8027;
  assign T_8032 = T_6928[27];
  assign T_8036 = ~ T_8032;
  assign T_8038 = T_8036 == 1'h0;
  assign T_8052 = T_3205_bits_data[27];
  assign GEN_3566 = {{27'd0}, pending_27};
  assign T_8067 = GEN_3566 << 27;
  assign GEN_3567 = {{1'd0}, T_8031};
  assign T_8071 = GEN_3567 | T_8067;
  assign T_8072 = T_6928[28];
  assign T_8076 = ~ T_8072;
  assign T_8078 = T_8076 == 1'h0;
  assign T_8092 = T_3205_bits_data[28];
  assign GEN_3568 = {{28'd0}, pending_28};
  assign T_8107 = GEN_3568 << 28;
  assign GEN_3569 = {{1'd0}, T_8071};
  assign T_8111 = GEN_3569 | T_8107;
  assign T_8112 = T_6928[29];
  assign T_8116 = ~ T_8112;
  assign T_8118 = T_8116 == 1'h0;
  assign T_8132 = T_3205_bits_data[29];
  assign GEN_3570 = {{29'd0}, pending_29};
  assign T_8147 = GEN_3570 << 29;
  assign GEN_3571 = {{1'd0}, T_8111};
  assign T_8151 = GEN_3571 | T_8147;
  assign T_8152 = T_6928[30];
  assign T_8156 = ~ T_8152;
  assign T_8158 = T_8156 == 1'h0;
  assign T_8172 = T_3205_bits_data[30];
  assign GEN_3572 = {{30'd0}, pending_30};
  assign T_8187 = GEN_3572 << 30;
  assign GEN_3573 = {{1'd0}, T_8151};
  assign T_8191 = GEN_3573 | T_8187;
  assign T_8192 = T_6928[31];
  assign T_8196 = ~ T_8192;
  assign T_8198 = T_8196 == 1'h0;
  assign T_8212 = T_3205_bits_data[31];
  assign GEN_3574 = {{31'd0}, pending_31};
  assign T_8227 = GEN_3574 << 31;
  assign GEN_3575 = {{1'd0}, T_8191};
  assign T_8231 = GEN_3575 | T_8227;
  assign T_8234 = T_6928 != 32'h0;
  assign T_8236 = ~ T_6928;
  assign T_8238 = T_8236 == 32'h0;
  assign T_8270 = {{29'd0}, priority_0};
  assign T_8291 = T_4344_33 & T_8238;
  assign GEN_61 = T_8291 ? T_3205_bits_data : {{29'd0}, priority_5};
  assign T_8310 = {{29'd0}, priority_5};
  assign T_8331 = T_4344_34 & T_8238;
  assign GEN_62 = T_8331 ? T_3205_bits_data : {{29'd0}, priority_10};
  assign T_8350 = {{29'd0}, priority_10};
  assign T_8371 = T_4344_35 & T_8238;
  assign GEN_63 = T_8371 ? T_3205_bits_data : {{29'd0}, priority_42};
  assign T_8390 = {{29'd0}, priority_42};
  assign T_8411 = T_4344_36 & T_8238;
  assign GEN_64 = T_8411 ? T_3205_bits_data : {{29'd0}, priority_24};
  assign T_8430 = {{29'd0}, priority_24};
  assign T_8451 = T_4344_37 & T_8238;
  assign GEN_65 = T_8451 ? T_3205_bits_data : {{29'd0}, priority_37};
  assign T_8470 = {{29'd0}, priority_37};
  assign T_8491 = T_4344_38 & T_8238;
  assign GEN_66 = T_8491 ? T_3205_bits_data : {{29'd0}, priority_25};
  assign T_8510 = {{29'd0}, priority_25};
  assign T_8531 = T_4344_39 & T_8238;
  assign GEN_67 = T_8531 ? T_3205_bits_data : {{29'd0}, priority_14};
  assign T_8550 = {{29'd0}, priority_14};
  assign T_8571 = T_4344_40 & T_8238;
  assign GEN_68 = T_8571 ? T_3205_bits_data : {{29'd0}, priority_20};
  assign T_8590 = {{29'd0}, priority_20};
  assign T_8611 = T_4344_41 & T_6958;
  assign GEN_69 = T_8611 ? T_6972 : enables_0_32;
  assign T_8651 = T_4344_42 & T_6998;
  assign GEN_70 = T_8651 ? T_7012 : enables_0_33;
  assign GEN_3576 = {{1'd0}, enables_0_33};
  assign T_8667 = GEN_3576 << 1;
  assign GEN_3577 = {{1'd0}, enables_0_32};
  assign T_8671 = GEN_3577 | T_8667;
  assign T_8691 = T_4344_43 & T_7038;
  assign GEN_71 = T_8691 ? T_7052 : enables_0_34;
  assign GEN_3578 = {{2'd0}, enables_0_34};
  assign T_8707 = GEN_3578 << 2;
  assign GEN_3579 = {{1'd0}, T_8671};
  assign T_8711 = GEN_3579 | T_8707;
  assign T_8731 = T_4344_44 & T_7078;
  assign GEN_72 = T_8731 ? T_7092 : enables_0_35;
  assign GEN_3580 = {{3'd0}, enables_0_35};
  assign T_8747 = GEN_3580 << 3;
  assign GEN_3581 = {{1'd0}, T_8711};
  assign T_8751 = GEN_3581 | T_8747;
  assign T_8771 = T_4344_45 & T_7118;
  assign GEN_73 = T_8771 ? T_7132 : enables_0_36;
  assign GEN_3582 = {{4'd0}, enables_0_36};
  assign T_8787 = GEN_3582 << 4;
  assign GEN_3583 = {{1'd0}, T_8751};
  assign T_8791 = GEN_3583 | T_8787;
  assign T_8811 = T_4344_46 & T_7158;
  assign GEN_74 = T_8811 ? T_7172 : enables_0_37;
  assign GEN_3584 = {{5'd0}, enables_0_37};
  assign T_8827 = GEN_3584 << 5;
  assign GEN_3585 = {{1'd0}, T_8791};
  assign T_8831 = GEN_3585 | T_8827;
  assign T_8851 = T_4344_47 & T_7198;
  assign GEN_75 = T_8851 ? T_7212 : enables_0_38;
  assign GEN_3586 = {{6'd0}, enables_0_38};
  assign T_8867 = GEN_3586 << 6;
  assign GEN_3587 = {{1'd0}, T_8831};
  assign T_8871 = GEN_3587 | T_8867;
  assign T_8891 = T_4344_48 & T_7238;
  assign GEN_76 = T_8891 ? T_7252 : enables_0_39;
  assign GEN_3588 = {{7'd0}, enables_0_39};
  assign T_8907 = GEN_3588 << 7;
  assign GEN_3589 = {{1'd0}, T_8871};
  assign T_8911 = GEN_3589 | T_8907;
  assign T_8931 = T_4344_49 & T_7278;
  assign GEN_77 = T_8931 ? T_7292 : enables_0_40;
  assign GEN_3590 = {{8'd0}, enables_0_40};
  assign T_8947 = GEN_3590 << 8;
  assign GEN_3591 = {{1'd0}, T_8911};
  assign T_8951 = GEN_3591 | T_8947;
  assign T_8971 = T_4344_50 & T_7318;
  assign GEN_78 = T_8971 ? T_7332 : enables_0_41;
  assign GEN_3592 = {{9'd0}, enables_0_41};
  assign T_8987 = GEN_3592 << 9;
  assign GEN_3593 = {{1'd0}, T_8951};
  assign T_8991 = GEN_3593 | T_8987;
  assign T_9011 = T_4344_51 & T_7358;
  assign GEN_79 = T_9011 ? T_7372 : enables_0_42;
  assign GEN_3594 = {{10'd0}, enables_0_42};
  assign T_9027 = GEN_3594 << 10;
  assign GEN_3595 = {{1'd0}, T_8991};
  assign T_9031 = GEN_3595 | T_9027;
  assign T_9051 = T_4344_52 & T_7398;
  assign GEN_80 = T_9051 ? T_7412 : enables_0_43;
  assign GEN_3596 = {{11'd0}, enables_0_43};
  assign T_9067 = GEN_3596 << 11;
  assign GEN_3597 = {{1'd0}, T_9031};
  assign T_9071 = GEN_3597 | T_9067;
  assign T_9091 = T_4344_53 & T_7438;
  assign GEN_81 = T_9091 ? T_7452 : enables_0_44;
  assign GEN_3598 = {{12'd0}, enables_0_44};
  assign T_9107 = GEN_3598 << 12;
  assign GEN_3599 = {{1'd0}, T_9071};
  assign T_9111 = GEN_3599 | T_9107;
  assign T_9131 = T_4344_54 & T_7478;
  assign GEN_82 = T_9131 ? T_7492 : enables_0_45;
  assign GEN_3600 = {{13'd0}, enables_0_45};
  assign T_9147 = GEN_3600 << 13;
  assign GEN_3601 = {{1'd0}, T_9111};
  assign T_9151 = GEN_3601 | T_9147;
  assign T_9171 = T_4344_55 & T_7518;
  assign GEN_83 = T_9171 ? T_7532 : enables_0_46;
  assign GEN_3602 = {{14'd0}, enables_0_46};
  assign T_9187 = GEN_3602 << 14;
  assign GEN_3603 = {{1'd0}, T_9151};
  assign T_9191 = GEN_3603 | T_9187;
  assign T_9211 = T_4344_56 & T_7558;
  assign GEN_84 = T_9211 ? T_7572 : enables_0_47;
  assign GEN_3604 = {{15'd0}, enables_0_47};
  assign T_9227 = GEN_3604 << 15;
  assign GEN_3605 = {{1'd0}, T_9191};
  assign T_9231 = GEN_3605 | T_9227;
  assign T_9251 = T_4344_57 & T_7598;
  assign GEN_85 = T_9251 ? T_7612 : enables_0_48;
  assign GEN_3606 = {{16'd0}, enables_0_48};
  assign T_9267 = GEN_3606 << 16;
  assign GEN_3607 = {{1'd0}, T_9231};
  assign T_9271 = GEN_3607 | T_9267;
  assign T_9291 = T_4344_58 & T_7638;
  assign GEN_86 = T_9291 ? T_7652 : enables_0_49;
  assign GEN_3608 = {{17'd0}, enables_0_49};
  assign T_9307 = GEN_3608 << 17;
  assign GEN_3609 = {{1'd0}, T_9271};
  assign T_9311 = GEN_3609 | T_9307;
  assign T_9331 = T_4344_59 & T_7678;
  assign GEN_87 = T_9331 ? T_7692 : enables_0_50;
  assign GEN_3610 = {{18'd0}, enables_0_50};
  assign T_9347 = GEN_3610 << 18;
  assign GEN_3611 = {{1'd0}, T_9311};
  assign T_9351 = GEN_3611 | T_9347;
  assign T_9371 = T_4344_60 & T_7718;
  assign GEN_88 = T_9371 ? T_7732 : enables_0_51;
  assign GEN_3612 = {{19'd0}, enables_0_51};
  assign T_9387 = GEN_3612 << 19;
  assign GEN_3613 = {{1'd0}, T_9351};
  assign T_9391 = GEN_3613 | T_9387;
  assign T_9411 = T_4344_61 & T_8238;
  assign GEN_89 = T_9411 ? T_3205_bits_data : {{29'd0}, priority_46};
  assign T_9430 = {{29'd0}, priority_46};
  assign T_9451 = T_4344_62 & T_8238;
  assign GEN_90 = T_9451 ? T_3205_bits_data : {{29'd0}, priority_29};
  assign T_9470 = {{29'd0}, priority_29};
  assign T_9487 = T_4339_63 & T_8234;
  assign GEN_0 = 1'h0;
  assign GEN_92 = 6'h1 == maxDevs_0 ? GEN_0 : GEN_9;
  assign GEN_93 = 6'h2 == maxDevs_0 ? GEN_0 : GEN_10;
  assign GEN_94 = 6'h3 == maxDevs_0 ? GEN_0 : GEN_11;
  assign GEN_95 = 6'h4 == maxDevs_0 ? GEN_0 : GEN_12;
  assign GEN_96 = 6'h5 == maxDevs_0 ? GEN_0 : GEN_13;
  assign GEN_97 = 6'h6 == maxDevs_0 ? GEN_0 : GEN_14;
  assign GEN_98 = 6'h7 == maxDevs_0 ? GEN_0 : GEN_15;
  assign GEN_99 = 6'h8 == maxDevs_0 ? GEN_0 : GEN_16;
  assign GEN_100 = 6'h9 == maxDevs_0 ? GEN_0 : GEN_17;
  assign GEN_101 = 6'ha == maxDevs_0 ? GEN_0 : GEN_18;
  assign GEN_102 = 6'hb == maxDevs_0 ? GEN_0 : GEN_19;
  assign GEN_103 = 6'hc == maxDevs_0 ? GEN_0 : GEN_20;
  assign GEN_104 = 6'hd == maxDevs_0 ? GEN_0 : GEN_21;
  assign GEN_105 = 6'he == maxDevs_0 ? GEN_0 : GEN_22;
  assign GEN_106 = 6'hf == maxDevs_0 ? GEN_0 : GEN_23;
  assign GEN_107 = 6'h10 == maxDevs_0 ? GEN_0 : GEN_24;
  assign GEN_108 = 6'h11 == maxDevs_0 ? GEN_0 : GEN_25;
  assign GEN_109 = 6'h12 == maxDevs_0 ? GEN_0 : GEN_26;
  assign GEN_110 = 6'h13 == maxDevs_0 ? GEN_0 : GEN_27;
  assign GEN_111 = 6'h14 == maxDevs_0 ? GEN_0 : GEN_28;
  assign GEN_112 = 6'h15 == maxDevs_0 ? GEN_0 : GEN_29;
  assign GEN_113 = 6'h16 == maxDevs_0 ? GEN_0 : GEN_30;
  assign GEN_114 = 6'h17 == maxDevs_0 ? GEN_0 : GEN_31;
  assign GEN_115 = 6'h18 == maxDevs_0 ? GEN_0 : GEN_32;
  assign GEN_116 = 6'h19 == maxDevs_0 ? GEN_0 : GEN_33;
  assign GEN_117 = 6'h1a == maxDevs_0 ? GEN_0 : GEN_34;
  assign GEN_118 = 6'h1b == maxDevs_0 ? GEN_0 : GEN_35;
  assign GEN_119 = 6'h1c == maxDevs_0 ? GEN_0 : GEN_36;
  assign GEN_120 = 6'h1d == maxDevs_0 ? GEN_0 : GEN_37;
  assign GEN_121 = 6'h1e == maxDevs_0 ? GEN_0 : GEN_38;
  assign GEN_122 = 6'h1f == maxDevs_0 ? GEN_0 : GEN_39;
  assign GEN_123 = 6'h20 == maxDevs_0 ? GEN_0 : GEN_40;
  assign GEN_124 = 6'h21 == maxDevs_0 ? GEN_0 : GEN_41;
  assign GEN_125 = 6'h22 == maxDevs_0 ? GEN_0 : GEN_42;
  assign GEN_126 = 6'h23 == maxDevs_0 ? GEN_0 : GEN_43;
  assign GEN_127 = 6'h24 == maxDevs_0 ? GEN_0 : GEN_44;
  assign GEN_128 = 6'h25 == maxDevs_0 ? GEN_0 : GEN_45;
  assign GEN_129 = 6'h26 == maxDevs_0 ? GEN_0 : GEN_46;
  assign GEN_130 = 6'h27 == maxDevs_0 ? GEN_0 : GEN_47;
  assign GEN_131 = 6'h28 == maxDevs_0 ? GEN_0 : GEN_48;
  assign GEN_132 = 6'h29 == maxDevs_0 ? GEN_0 : GEN_49;
  assign GEN_133 = 6'h2a == maxDevs_0 ? GEN_0 : GEN_50;
  assign GEN_134 = 6'h2b == maxDevs_0 ? GEN_0 : GEN_51;
  assign GEN_135 = 6'h2c == maxDevs_0 ? GEN_0 : GEN_52;
  assign GEN_136 = 6'h2d == maxDevs_0 ? GEN_0 : GEN_53;
  assign GEN_137 = 6'h2e == maxDevs_0 ? GEN_0 : GEN_54;
  assign GEN_138 = 6'h2f == maxDevs_0 ? GEN_0 : GEN_55;
  assign GEN_139 = 6'h30 == maxDevs_0 ? GEN_0 : GEN_56;
  assign GEN_140 = 6'h31 == maxDevs_0 ? GEN_0 : GEN_57;
  assign GEN_141 = 6'h32 == maxDevs_0 ? GEN_0 : GEN_58;
  assign GEN_142 = 6'h33 == maxDevs_0 ? GEN_0 : GEN_59;
  assign GEN_144 = T_9487 ? GEN_92 : GEN_9;
  assign GEN_145 = T_9487 ? GEN_93 : GEN_10;
  assign GEN_146 = T_9487 ? GEN_94 : GEN_11;
  assign GEN_147 = T_9487 ? GEN_95 : GEN_12;
  assign GEN_148 = T_9487 ? GEN_96 : GEN_13;
  assign GEN_149 = T_9487 ? GEN_97 : GEN_14;
  assign GEN_150 = T_9487 ? GEN_98 : GEN_15;
  assign GEN_151 = T_9487 ? GEN_99 : GEN_16;
  assign GEN_152 = T_9487 ? GEN_100 : GEN_17;
  assign GEN_153 = T_9487 ? GEN_101 : GEN_18;
  assign GEN_154 = T_9487 ? GEN_102 : GEN_19;
  assign GEN_155 = T_9487 ? GEN_103 : GEN_20;
  assign GEN_156 = T_9487 ? GEN_104 : GEN_21;
  assign GEN_157 = T_9487 ? GEN_105 : GEN_22;
  assign GEN_158 = T_9487 ? GEN_106 : GEN_23;
  assign GEN_159 = T_9487 ? GEN_107 : GEN_24;
  assign GEN_160 = T_9487 ? GEN_108 : GEN_25;
  assign GEN_161 = T_9487 ? GEN_109 : GEN_26;
  assign GEN_162 = T_9487 ? GEN_110 : GEN_27;
  assign GEN_163 = T_9487 ? GEN_111 : GEN_28;
  assign GEN_164 = T_9487 ? GEN_112 : GEN_29;
  assign GEN_165 = T_9487 ? GEN_113 : GEN_30;
  assign GEN_166 = T_9487 ? GEN_114 : GEN_31;
  assign GEN_167 = T_9487 ? GEN_115 : GEN_32;
  assign GEN_168 = T_9487 ? GEN_116 : GEN_33;
  assign GEN_169 = T_9487 ? GEN_117 : GEN_34;
  assign GEN_170 = T_9487 ? GEN_118 : GEN_35;
  assign GEN_171 = T_9487 ? GEN_119 : GEN_36;
  assign GEN_172 = T_9487 ? GEN_120 : GEN_37;
  assign GEN_173 = T_9487 ? GEN_121 : GEN_38;
  assign GEN_174 = T_9487 ? GEN_122 : GEN_39;
  assign GEN_175 = T_9487 ? GEN_123 : GEN_40;
  assign GEN_176 = T_9487 ? GEN_124 : GEN_41;
  assign GEN_177 = T_9487 ? GEN_125 : GEN_42;
  assign GEN_178 = T_9487 ? GEN_126 : GEN_43;
  assign GEN_179 = T_9487 ? GEN_127 : GEN_44;
  assign GEN_180 = T_9487 ? GEN_128 : GEN_45;
  assign GEN_181 = T_9487 ? GEN_129 : GEN_46;
  assign GEN_182 = T_9487 ? GEN_130 : GEN_47;
  assign GEN_183 = T_9487 ? GEN_131 : GEN_48;
  assign GEN_184 = T_9487 ? GEN_132 : GEN_49;
  assign GEN_185 = T_9487 ? GEN_133 : GEN_50;
  assign GEN_186 = T_9487 ? GEN_134 : GEN_51;
  assign GEN_187 = T_9487 ? GEN_135 : GEN_52;
  assign GEN_188 = T_9487 ? GEN_136 : GEN_53;
  assign GEN_189 = T_9487 ? GEN_137 : GEN_54;
  assign GEN_190 = T_9487 ? GEN_138 : GEN_55;
  assign GEN_191 = T_9487 ? GEN_139 : GEN_56;
  assign GEN_192 = T_9487 ? GEN_140 : GEN_57;
  assign GEN_193 = T_9487 ? GEN_141 : GEN_58;
  assign GEN_194 = T_9487 ? GEN_142 : GEN_59;
  assign GEN_195 = T_9487 ? 6'h0 : T_3102;
  assign T_9494 = T_4344_63 & T_8238;
  assign T_9497 = T_3205_bits_data[5:0];
  assign GEN_1 = GEN_246;
  assign GEN_196 = 6'h1 == T_9497 ? enables_0_1 : enables_0_0;
  assign GEN_197 = 6'h2 == T_9497 ? enables_0_2 : GEN_196;
  assign GEN_198 = 6'h3 == T_9497 ? enables_0_3 : GEN_197;
  assign GEN_199 = 6'h4 == T_9497 ? enables_0_4 : GEN_198;
  assign GEN_200 = 6'h5 == T_9497 ? enables_0_5 : GEN_199;
  assign GEN_201 = 6'h6 == T_9497 ? enables_0_6 : GEN_200;
  assign GEN_202 = 6'h7 == T_9497 ? enables_0_7 : GEN_201;
  assign GEN_203 = 6'h8 == T_9497 ? enables_0_8 : GEN_202;
  assign GEN_204 = 6'h9 == T_9497 ? enables_0_9 : GEN_203;
  assign GEN_205 = 6'ha == T_9497 ? enables_0_10 : GEN_204;
  assign GEN_206 = 6'hb == T_9497 ? enables_0_11 : GEN_205;
  assign GEN_207 = 6'hc == T_9497 ? enables_0_12 : GEN_206;
  assign GEN_208 = 6'hd == T_9497 ? enables_0_13 : GEN_207;
  assign GEN_209 = 6'he == T_9497 ? enables_0_14 : GEN_208;
  assign GEN_210 = 6'hf == T_9497 ? enables_0_15 : GEN_209;
  assign GEN_211 = 6'h10 == T_9497 ? enables_0_16 : GEN_210;
  assign GEN_212 = 6'h11 == T_9497 ? enables_0_17 : GEN_211;
  assign GEN_213 = 6'h12 == T_9497 ? enables_0_18 : GEN_212;
  assign GEN_214 = 6'h13 == T_9497 ? enables_0_19 : GEN_213;
  assign GEN_215 = 6'h14 == T_9497 ? enables_0_20 : GEN_214;
  assign GEN_216 = 6'h15 == T_9497 ? enables_0_21 : GEN_215;
  assign GEN_217 = 6'h16 == T_9497 ? enables_0_22 : GEN_216;
  assign GEN_218 = 6'h17 == T_9497 ? enables_0_23 : GEN_217;
  assign GEN_219 = 6'h18 == T_9497 ? enables_0_24 : GEN_218;
  assign GEN_220 = 6'h19 == T_9497 ? enables_0_25 : GEN_219;
  assign GEN_221 = 6'h1a == T_9497 ? enables_0_26 : GEN_220;
  assign GEN_222 = 6'h1b == T_9497 ? enables_0_27 : GEN_221;
  assign GEN_223 = 6'h1c == T_9497 ? enables_0_28 : GEN_222;
  assign GEN_224 = 6'h1d == T_9497 ? enables_0_29 : GEN_223;
  assign GEN_225 = 6'h1e == T_9497 ? enables_0_30 : GEN_224;
  assign GEN_226 = 6'h1f == T_9497 ? enables_0_31 : GEN_225;
  assign GEN_227 = 6'h20 == T_9497 ? enables_0_32 : GEN_226;
  assign GEN_228 = 6'h21 == T_9497 ? enables_0_33 : GEN_227;
  assign GEN_229 = 6'h22 == T_9497 ? enables_0_34 : GEN_228;
  assign GEN_230 = 6'h23 == T_9497 ? enables_0_35 : GEN_229;
  assign GEN_231 = 6'h24 == T_9497 ? enables_0_36 : GEN_230;
  assign GEN_232 = 6'h25 == T_9497 ? enables_0_37 : GEN_231;
  assign GEN_233 = 6'h26 == T_9497 ? enables_0_38 : GEN_232;
  assign GEN_234 = 6'h27 == T_9497 ? enables_0_39 : GEN_233;
  assign GEN_235 = 6'h28 == T_9497 ? enables_0_40 : GEN_234;
  assign GEN_236 = 6'h29 == T_9497 ? enables_0_41 : GEN_235;
  assign GEN_237 = 6'h2a == T_9497 ? enables_0_42 : GEN_236;
  assign GEN_238 = 6'h2b == T_9497 ? enables_0_43 : GEN_237;
  assign GEN_239 = 6'h2c == T_9497 ? enables_0_44 : GEN_238;
  assign GEN_240 = 6'h2d == T_9497 ? enables_0_45 : GEN_239;
  assign GEN_241 = 6'h2e == T_9497 ? enables_0_46 : GEN_240;
  assign GEN_242 = 6'h2f == T_9497 ? enables_0_47 : GEN_241;
  assign GEN_243 = 6'h30 == T_9497 ? enables_0_48 : GEN_242;
  assign GEN_244 = 6'h31 == T_9497 ? enables_0_49 : GEN_243;
  assign GEN_245 = 6'h32 == T_9497 ? enables_0_50 : GEN_244;
  assign GEN_246 = 6'h33 == T_9497 ? enables_0_51 : GEN_245;
  assign T_9498 = T_9494 & GEN_1;
  assign T_9500 = T_3205_bits_data - 32'h1;
  assign T_9501 = T_9500[31:0];
  assign T_9515 = T_9501[5:0];
  assign GEN_2 = 1'h1;
  assign GEN_247 = 6'h0 == T_9515 ? GEN_2 : 1'h0;
  assign GEN_248 = 6'h1 == T_9515 ? GEN_2 : 1'h0;
  assign GEN_249 = 6'h2 == T_9515 ? GEN_2 : 1'h0;
  assign GEN_250 = 6'h3 == T_9515 ? GEN_2 : 1'h0;
  assign GEN_251 = 6'h4 == T_9515 ? GEN_2 : 1'h0;
  assign GEN_252 = 6'h5 == T_9515 ? GEN_2 : 1'h0;
  assign GEN_253 = 6'h6 == T_9515 ? GEN_2 : 1'h0;
  assign GEN_254 = 6'h7 == T_9515 ? GEN_2 : 1'h0;
  assign GEN_255 = 6'h8 == T_9515 ? GEN_2 : 1'h0;
  assign GEN_256 = 6'h9 == T_9515 ? GEN_2 : 1'h0;
  assign GEN_257 = 6'ha == T_9515 ? GEN_2 : 1'h0;
  assign GEN_258 = 6'hb == T_9515 ? GEN_2 : 1'h0;
  assign GEN_259 = 6'hc == T_9515 ? GEN_2 : 1'h0;
  assign GEN_260 = 6'hd == T_9515 ? GEN_2 : 1'h0;
  assign GEN_261 = 6'he == T_9515 ? GEN_2 : 1'h0;
  assign GEN_262 = 6'hf == T_9515 ? GEN_2 : 1'h0;
  assign GEN_263 = 6'h10 == T_9515 ? GEN_2 : 1'h0;
  assign GEN_264 = 6'h11 == T_9515 ? GEN_2 : 1'h0;
  assign GEN_265 = 6'h12 == T_9515 ? GEN_2 : 1'h0;
  assign GEN_266 = 6'h13 == T_9515 ? GEN_2 : 1'h0;
  assign GEN_267 = 6'h14 == T_9515 ? GEN_2 : 1'h0;
  assign GEN_268 = 6'h15 == T_9515 ? GEN_2 : 1'h0;
  assign GEN_269 = 6'h16 == T_9515 ? GEN_2 : 1'h0;
  assign GEN_270 = 6'h17 == T_9515 ? GEN_2 : 1'h0;
  assign GEN_271 = 6'h18 == T_9515 ? GEN_2 : 1'h0;
  assign GEN_272 = 6'h19 == T_9515 ? GEN_2 : 1'h0;
  assign GEN_273 = 6'h1a == T_9515 ? GEN_2 : 1'h0;
  assign GEN_274 = 6'h1b == T_9515 ? GEN_2 : 1'h0;
  assign GEN_275 = 6'h1c == T_9515 ? GEN_2 : 1'h0;
  assign GEN_276 = 6'h1d == T_9515 ? GEN_2 : 1'h0;
  assign GEN_277 = 6'h1e == T_9515 ? GEN_2 : 1'h0;
  assign GEN_278 = 6'h1f == T_9515 ? GEN_2 : 1'h0;
  assign GEN_279 = 6'h20 == T_9515 ? GEN_2 : 1'h0;
  assign GEN_280 = 6'h21 == T_9515 ? GEN_2 : 1'h0;
  assign GEN_281 = 6'h22 == T_9515 ? GEN_2 : 1'h0;
  assign GEN_282 = 6'h23 == T_9515 ? GEN_2 : 1'h0;
  assign GEN_283 = 6'h24 == T_9515 ? GEN_2 : 1'h0;
  assign GEN_284 = 6'h25 == T_9515 ? GEN_2 : 1'h0;
  assign GEN_285 = 6'h26 == T_9515 ? GEN_2 : 1'h0;
  assign GEN_286 = 6'h27 == T_9515 ? GEN_2 : 1'h0;
  assign GEN_287 = 6'h28 == T_9515 ? GEN_2 : 1'h0;
  assign GEN_288 = 6'h29 == T_9515 ? GEN_2 : 1'h0;
  assign GEN_289 = 6'h2a == T_9515 ? GEN_2 : 1'h0;
  assign GEN_290 = 6'h2b == T_9515 ? GEN_2 : 1'h0;
  assign GEN_291 = 6'h2c == T_9515 ? GEN_2 : 1'h0;
  assign GEN_292 = 6'h2d == T_9515 ? GEN_2 : 1'h0;
  assign GEN_293 = 6'h2e == T_9515 ? GEN_2 : 1'h0;
  assign GEN_294 = 6'h2f == T_9515 ? GEN_2 : 1'h0;
  assign GEN_295 = 6'h30 == T_9515 ? GEN_2 : 1'h0;
  assign GEN_296 = 6'h31 == T_9515 ? GEN_2 : 1'h0;
  assign GEN_297 = 6'h32 == T_9515 ? GEN_2 : 1'h0;
  assign GEN_298 = T_9498 ? GEN_247 : 1'h0;
  assign GEN_299 = T_9498 ? GEN_248 : 1'h0;
  assign GEN_300 = T_9498 ? GEN_249 : 1'h0;
  assign GEN_301 = T_9498 ? GEN_250 : 1'h0;
  assign GEN_302 = T_9498 ? GEN_251 : 1'h0;
  assign GEN_303 = T_9498 ? GEN_252 : 1'h0;
  assign GEN_304 = T_9498 ? GEN_253 : 1'h0;
  assign GEN_305 = T_9498 ? GEN_254 : 1'h0;
  assign GEN_306 = T_9498 ? GEN_255 : 1'h0;
  assign GEN_307 = T_9498 ? GEN_256 : 1'h0;
  assign GEN_308 = T_9498 ? GEN_257 : 1'h0;
  assign GEN_309 = T_9498 ? GEN_258 : 1'h0;
  assign GEN_310 = T_9498 ? GEN_259 : 1'h0;
  assign GEN_311 = T_9498 ? GEN_260 : 1'h0;
  assign GEN_312 = T_9498 ? GEN_261 : 1'h0;
  assign GEN_313 = T_9498 ? GEN_262 : 1'h0;
  assign GEN_314 = T_9498 ? GEN_263 : 1'h0;
  assign GEN_315 = T_9498 ? GEN_264 : 1'h0;
  assign GEN_316 = T_9498 ? GEN_265 : 1'h0;
  assign GEN_317 = T_9498 ? GEN_266 : 1'h0;
  assign GEN_318 = T_9498 ? GEN_267 : 1'h0;
  assign GEN_319 = T_9498 ? GEN_268 : 1'h0;
  assign GEN_320 = T_9498 ? GEN_269 : 1'h0;
  assign GEN_321 = T_9498 ? GEN_270 : 1'h0;
  assign GEN_322 = T_9498 ? GEN_271 : 1'h0;
  assign GEN_323 = T_9498 ? GEN_272 : 1'h0;
  assign GEN_324 = T_9498 ? GEN_273 : 1'h0;
  assign GEN_325 = T_9498 ? GEN_274 : 1'h0;
  assign GEN_326 = T_9498 ? GEN_275 : 1'h0;
  assign GEN_327 = T_9498 ? GEN_276 : 1'h0;
  assign GEN_328 = T_9498 ? GEN_277 : 1'h0;
  assign GEN_329 = T_9498 ? GEN_278 : 1'h0;
  assign GEN_330 = T_9498 ? GEN_279 : 1'h0;
  assign GEN_331 = T_9498 ? GEN_280 : 1'h0;
  assign GEN_332 = T_9498 ? GEN_281 : 1'h0;
  assign GEN_333 = T_9498 ? GEN_282 : 1'h0;
  assign GEN_334 = T_9498 ? GEN_283 : 1'h0;
  assign GEN_335 = T_9498 ? GEN_284 : 1'h0;
  assign GEN_336 = T_9498 ? GEN_285 : 1'h0;
  assign GEN_337 = T_9498 ? GEN_286 : 1'h0;
  assign GEN_338 = T_9498 ? GEN_287 : 1'h0;
  assign GEN_339 = T_9498 ? GEN_288 : 1'h0;
  assign GEN_340 = T_9498 ? GEN_289 : 1'h0;
  assign GEN_341 = T_9498 ? GEN_290 : 1'h0;
  assign GEN_342 = T_9498 ? GEN_291 : 1'h0;
  assign GEN_343 = T_9498 ? GEN_292 : 1'h0;
  assign GEN_344 = T_9498 ? GEN_293 : 1'h0;
  assign GEN_345 = T_9498 ? GEN_294 : 1'h0;
  assign GEN_346 = T_9498 ? GEN_295 : 1'h0;
  assign GEN_347 = T_9498 ? GEN_296 : 1'h0;
  assign GEN_348 = T_9498 ? GEN_297 : 1'h0;
  assign T_9533 = {{26'd0}, maxDevs_0};
  assign T_9554 = T_4344_64 & T_8238;
  assign GEN_349 = T_9554 ? T_3205_bits_data : {{29'd0}, priority_1};
  assign T_9573 = {{29'd0}, priority_1};
  assign T_9594 = T_4344_65 & T_8238;
  assign GEN_350 = T_9594 ? T_3205_bits_data : {{29'd0}, priority_6};
  assign T_9613 = {{29'd0}, priority_6};
  assign T_9634 = T_4344_66 & T_8238;
  assign GEN_351 = T_9634 ? T_3205_bits_data : {{29'd0}, priority_28};
  assign T_9653 = {{29'd0}, priority_28};
  assign T_9674 = T_4344_67 & T_8238;
  assign GEN_352 = T_9674 ? T_3205_bits_data : {{29'd0}, priority_38};
  assign T_9693 = {{29'd0}, priority_38};
  assign T_9714 = T_4344_68 & T_8238;
  assign GEN_353 = T_9714 ? T_3205_bits_data : {{29'd0}, priority_21};
  assign T_9733 = {{29'd0}, priority_21};
  assign T_9754 = T_4344_69 & T_8238;
  assign GEN_354 = T_9754 ? T_3205_bits_data : {{29'd0}, priority_33};
  assign T_9773 = {{29'd0}, priority_33};
  assign T_9794 = T_4344_70 & T_8238;
  assign GEN_355 = T_9794 ? T_3205_bits_data : {{29'd0}, priority_9};
  assign T_9813 = {{29'd0}, priority_9};
  assign T_9834 = T_4344_71 & T_8238;
  assign GEN_356 = T_9834 ? T_3205_bits_data : {{29'd0}, priority_13};
  assign T_9853 = {{29'd0}, priority_13};
  assign T_9874 = T_4344_72 & T_8238;
  assign GEN_357 = T_9874 ? T_3205_bits_data : {{29'd0}, priority_41};
  assign T_9893 = {{29'd0}, priority_41};
  assign T_9914 = T_4344_73 & T_8238;
  assign GEN_358 = T_9914 ? T_3205_bits_data : {{29'd0}, priority_2};
  assign T_9933 = {{29'd0}, priority_2};
  assign T_9954 = T_4344_74 & T_8238;
  assign GEN_359 = T_9954 ? T_3205_bits_data : {{29'd0}, priority_32};
  assign T_9973 = {{29'd0}, priority_32};
  assign T_9994 = T_4344_75 & T_8238;
  assign GEN_360 = T_9994 ? T_3205_bits_data : {{29'd0}, priority_34};
  assign T_10013 = {{29'd0}, priority_34};
  assign T_10034 = T_4344_76 & T_8238;
  assign GEN_361 = T_10034 ? T_3205_bits_data : {{29'd0}, priority_45};
  assign T_10053 = {{29'd0}, priority_45};
  assign T_10074 = T_4344_77 & T_8238;
  assign GEN_362 = T_10074 ? T_3205_bits_data : {{29'd0}, priority_17};
  assign T_10093 = {{29'd0}, priority_17};
  assign T_10114 = T_4344_78 & T_8238;
  assign GEN_363 = T_10114 ? T_3205_bits_data : {{29'd0}, threshold_0};
  assign T_10133 = {{29'd0}, threshold_0};
  assign T_10194 = T_4344_80 & T_6998;
  assign GEN_365 = T_10194 ? T_7012 : enables_0_1;
  assign GEN_3614 = {{1'd0}, enables_0_1};
  assign T_10210 = GEN_3614 << 1;
  assign GEN_3615 = {{1'd0}, enables_0_0};
  assign T_10214 = GEN_3615 | T_10210;
  assign T_10234 = T_4344_81 & T_7038;
  assign GEN_366 = T_10234 ? T_7052 : enables_0_2;
  assign GEN_3616 = {{2'd0}, enables_0_2};
  assign T_10250 = GEN_3616 << 2;
  assign GEN_3617 = {{1'd0}, T_10214};
  assign T_10254 = GEN_3617 | T_10250;
  assign T_10274 = T_4344_82 & T_7078;
  assign GEN_367 = T_10274 ? T_7092 : enables_0_3;
  assign GEN_3618 = {{3'd0}, enables_0_3};
  assign T_10290 = GEN_3618 << 3;
  assign GEN_3619 = {{1'd0}, T_10254};
  assign T_10294 = GEN_3619 | T_10290;
  assign T_10314 = T_4344_83 & T_7118;
  assign GEN_368 = T_10314 ? T_7132 : enables_0_4;
  assign GEN_3620 = {{4'd0}, enables_0_4};
  assign T_10330 = GEN_3620 << 4;
  assign GEN_3621 = {{1'd0}, T_10294};
  assign T_10334 = GEN_3621 | T_10330;
  assign T_10354 = T_4344_84 & T_7158;
  assign GEN_369 = T_10354 ? T_7172 : enables_0_5;
  assign GEN_3622 = {{5'd0}, enables_0_5};
  assign T_10370 = GEN_3622 << 5;
  assign GEN_3623 = {{1'd0}, T_10334};
  assign T_10374 = GEN_3623 | T_10370;
  assign T_10394 = T_4344_85 & T_7198;
  assign GEN_370 = T_10394 ? T_7212 : enables_0_6;
  assign GEN_3624 = {{6'd0}, enables_0_6};
  assign T_10410 = GEN_3624 << 6;
  assign GEN_3625 = {{1'd0}, T_10374};
  assign T_10414 = GEN_3625 | T_10410;
  assign T_10434 = T_4344_86 & T_7238;
  assign GEN_371 = T_10434 ? T_7252 : enables_0_7;
  assign GEN_3626 = {{7'd0}, enables_0_7};
  assign T_10450 = GEN_3626 << 7;
  assign GEN_3627 = {{1'd0}, T_10414};
  assign T_10454 = GEN_3627 | T_10450;
  assign T_10474 = T_4344_87 & T_7278;
  assign GEN_372 = T_10474 ? T_7292 : enables_0_8;
  assign GEN_3628 = {{8'd0}, enables_0_8};
  assign T_10490 = GEN_3628 << 8;
  assign GEN_3629 = {{1'd0}, T_10454};
  assign T_10494 = GEN_3629 | T_10490;
  assign T_10514 = T_4344_88 & T_7318;
  assign GEN_373 = T_10514 ? T_7332 : enables_0_9;
  assign GEN_3630 = {{9'd0}, enables_0_9};
  assign T_10530 = GEN_3630 << 9;
  assign GEN_3631 = {{1'd0}, T_10494};
  assign T_10534 = GEN_3631 | T_10530;
  assign T_10554 = T_4344_89 & T_7358;
  assign GEN_374 = T_10554 ? T_7372 : enables_0_10;
  assign GEN_3632 = {{10'd0}, enables_0_10};
  assign T_10570 = GEN_3632 << 10;
  assign GEN_3633 = {{1'd0}, T_10534};
  assign T_10574 = GEN_3633 | T_10570;
  assign T_10594 = T_4344_90 & T_7398;
  assign GEN_375 = T_10594 ? T_7412 : enables_0_11;
  assign GEN_3634 = {{11'd0}, enables_0_11};
  assign T_10610 = GEN_3634 << 11;
  assign GEN_3635 = {{1'd0}, T_10574};
  assign T_10614 = GEN_3635 | T_10610;
  assign T_10634 = T_4344_91 & T_7438;
  assign GEN_376 = T_10634 ? T_7452 : enables_0_12;
  assign GEN_3636 = {{12'd0}, enables_0_12};
  assign T_10650 = GEN_3636 << 12;
  assign GEN_3637 = {{1'd0}, T_10614};
  assign T_10654 = GEN_3637 | T_10650;
  assign T_10674 = T_4344_92 & T_7478;
  assign GEN_377 = T_10674 ? T_7492 : enables_0_13;
  assign GEN_3638 = {{13'd0}, enables_0_13};
  assign T_10690 = GEN_3638 << 13;
  assign GEN_3639 = {{1'd0}, T_10654};
  assign T_10694 = GEN_3639 | T_10690;
  assign T_10714 = T_4344_93 & T_7518;
  assign GEN_378 = T_10714 ? T_7532 : enables_0_14;
  assign GEN_3640 = {{14'd0}, enables_0_14};
  assign T_10730 = GEN_3640 << 14;
  assign GEN_3641 = {{1'd0}, T_10694};
  assign T_10734 = GEN_3641 | T_10730;
  assign T_10754 = T_4344_94 & T_7558;
  assign GEN_379 = T_10754 ? T_7572 : enables_0_15;
  assign GEN_3642 = {{15'd0}, enables_0_15};
  assign T_10770 = GEN_3642 << 15;
  assign GEN_3643 = {{1'd0}, T_10734};
  assign T_10774 = GEN_3643 | T_10770;
  assign T_10794 = T_4344_95 & T_7598;
  assign GEN_380 = T_10794 ? T_7612 : enables_0_16;
  assign GEN_3644 = {{16'd0}, enables_0_16};
  assign T_10810 = GEN_3644 << 16;
  assign GEN_3645 = {{1'd0}, T_10774};
  assign T_10814 = GEN_3645 | T_10810;
  assign T_10834 = T_4344_96 & T_7638;
  assign GEN_381 = T_10834 ? T_7652 : enables_0_17;
  assign GEN_3646 = {{17'd0}, enables_0_17};
  assign T_10850 = GEN_3646 << 17;
  assign GEN_3647 = {{1'd0}, T_10814};
  assign T_10854 = GEN_3647 | T_10850;
  assign T_10874 = T_4344_97 & T_7678;
  assign GEN_382 = T_10874 ? T_7692 : enables_0_18;
  assign GEN_3648 = {{18'd0}, enables_0_18};
  assign T_10890 = GEN_3648 << 18;
  assign GEN_3649 = {{1'd0}, T_10854};
  assign T_10894 = GEN_3649 | T_10890;
  assign T_10914 = T_4344_98 & T_7718;
  assign GEN_383 = T_10914 ? T_7732 : enables_0_19;
  assign GEN_3650 = {{19'd0}, enables_0_19};
  assign T_10930 = GEN_3650 << 19;
  assign GEN_3651 = {{1'd0}, T_10894};
  assign T_10934 = GEN_3651 | T_10930;
  assign T_10954 = T_4344_99 & T_7758;
  assign GEN_384 = T_10954 ? T_7772 : enables_0_20;
  assign GEN_3652 = {{20'd0}, enables_0_20};
  assign T_10970 = GEN_3652 << 20;
  assign GEN_3653 = {{1'd0}, T_10934};
  assign T_10974 = GEN_3653 | T_10970;
  assign T_10994 = T_4344_100 & T_7798;
  assign GEN_385 = T_10994 ? T_7812 : enables_0_21;
  assign GEN_3654 = {{21'd0}, enables_0_21};
  assign T_11010 = GEN_3654 << 21;
  assign GEN_3655 = {{1'd0}, T_10974};
  assign T_11014 = GEN_3655 | T_11010;
  assign T_11034 = T_4344_101 & T_7838;
  assign GEN_386 = T_11034 ? T_7852 : enables_0_22;
  assign GEN_3656 = {{22'd0}, enables_0_22};
  assign T_11050 = GEN_3656 << 22;
  assign GEN_3657 = {{1'd0}, T_11014};
  assign T_11054 = GEN_3657 | T_11050;
  assign T_11074 = T_4344_102 & T_7878;
  assign GEN_387 = T_11074 ? T_7892 : enables_0_23;
  assign GEN_3658 = {{23'd0}, enables_0_23};
  assign T_11090 = GEN_3658 << 23;
  assign GEN_3659 = {{1'd0}, T_11054};
  assign T_11094 = GEN_3659 | T_11090;
  assign T_11114 = T_4344_103 & T_7918;
  assign GEN_388 = T_11114 ? T_7932 : enables_0_24;
  assign GEN_3660 = {{24'd0}, enables_0_24};
  assign T_11130 = GEN_3660 << 24;
  assign GEN_3661 = {{1'd0}, T_11094};
  assign T_11134 = GEN_3661 | T_11130;
  assign T_11154 = T_4344_104 & T_7958;
  assign GEN_389 = T_11154 ? T_7972 : enables_0_25;
  assign GEN_3662 = {{25'd0}, enables_0_25};
  assign T_11170 = GEN_3662 << 25;
  assign GEN_3663 = {{1'd0}, T_11134};
  assign T_11174 = GEN_3663 | T_11170;
  assign T_11194 = T_4344_105 & T_7998;
  assign GEN_390 = T_11194 ? T_8012 : enables_0_26;
  assign GEN_3664 = {{26'd0}, enables_0_26};
  assign T_11210 = GEN_3664 << 26;
  assign GEN_3665 = {{1'd0}, T_11174};
  assign T_11214 = GEN_3665 | T_11210;
  assign T_11234 = T_4344_106 & T_8038;
  assign GEN_391 = T_11234 ? T_8052 : enables_0_27;
  assign GEN_3666 = {{27'd0}, enables_0_27};
  assign T_11250 = GEN_3666 << 27;
  assign GEN_3667 = {{1'd0}, T_11214};
  assign T_11254 = GEN_3667 | T_11250;
  assign T_11274 = T_4344_107 & T_8078;
  assign GEN_392 = T_11274 ? T_8092 : enables_0_28;
  assign GEN_3668 = {{28'd0}, enables_0_28};
  assign T_11290 = GEN_3668 << 28;
  assign GEN_3669 = {{1'd0}, T_11254};
  assign T_11294 = GEN_3669 | T_11290;
  assign T_11314 = T_4344_108 & T_8118;
  assign GEN_393 = T_11314 ? T_8132 : enables_0_29;
  assign GEN_3670 = {{29'd0}, enables_0_29};
  assign T_11330 = GEN_3670 << 29;
  assign GEN_3671 = {{1'd0}, T_11294};
  assign T_11334 = GEN_3671 | T_11330;
  assign T_11354 = T_4344_109 & T_8158;
  assign GEN_394 = T_11354 ? T_8172 : enables_0_30;
  assign GEN_3672 = {{30'd0}, enables_0_30};
  assign T_11370 = GEN_3672 << 30;
  assign GEN_3673 = {{1'd0}, T_11334};
  assign T_11374 = GEN_3673 | T_11370;
  assign T_11394 = T_4344_110 & T_8198;
  assign GEN_395 = T_11394 ? T_8212 : enables_0_31;
  assign GEN_3674 = {{31'd0}, enables_0_31};
  assign T_11410 = GEN_3674 << 31;
  assign GEN_3675 = {{1'd0}, T_11374};
  assign T_11414 = GEN_3675 | T_11410;
  assign T_11434 = T_4344_111 & T_8238;
  assign GEN_396 = T_11434 ? T_3205_bits_data : {{29'd0}, priority_22};
  assign T_11453 = {{29'd0}, priority_22};
  assign T_11474 = T_4344_112 & T_8238;
  assign GEN_397 = T_11474 ? T_3205_bits_data : {{29'd0}, priority_44};
  assign T_11493 = {{29'd0}, priority_44};
  assign T_11514 = T_4344_113 & T_8238;
  assign GEN_398 = T_11514 ? T_3205_bits_data : {{29'd0}, priority_27};
  assign T_11533 = {{29'd0}, priority_27};
  assign T_11554 = T_4344_114 & T_8238;
  assign GEN_399 = T_11554 ? T_3205_bits_data : {{29'd0}, priority_12};
  assign T_11573 = {{29'd0}, priority_12};
  assign T_11594 = T_4344_115 & T_8238;
  assign GEN_400 = T_11594 ? T_3205_bits_data : {{29'd0}, priority_49};
  assign T_11613 = {{29'd0}, priority_49};
  assign T_11634 = T_4344_116 & T_8238;
  assign GEN_401 = T_11634 ? T_3205_bits_data : {{29'd0}, priority_7};
  assign T_11653 = {{29'd0}, priority_7};
  assign T_11674 = T_4344_117 & T_8238;
  assign GEN_402 = T_11674 ? T_3205_bits_data : {{29'd0}, priority_39};
  assign T_11693 = {{29'd0}, priority_39};
  assign T_11714 = T_4344_118 & T_8238;
  assign GEN_403 = T_11714 ? T_3205_bits_data : {{29'd0}, priority_3};
  assign T_11733 = {{29'd0}, priority_3};
  assign T_11754 = T_4344_119 & T_8238;
  assign GEN_404 = T_11754 ? T_3205_bits_data : {{29'd0}, priority_35};
  assign T_11773 = {{29'd0}, priority_35};
  assign T_11794 = T_4344_120 & T_8238;
  assign GEN_405 = T_11794 ? T_3205_bits_data : {{29'd0}, priority_48};
  assign T_11813 = {{29'd0}, priority_48};
  assign GEN_3676 = {{1'd0}, pending_33};
  assign T_11890 = GEN_3676 << 1;
  assign GEN_3677 = {{1'd0}, pending_32};
  assign T_11894 = GEN_3677 | T_11890;
  assign GEN_3678 = {{2'd0}, pending_34};
  assign T_11930 = GEN_3678 << 2;
  assign GEN_3679 = {{1'd0}, T_11894};
  assign T_11934 = GEN_3679 | T_11930;
  assign GEN_3680 = {{3'd0}, pending_35};
  assign T_11970 = GEN_3680 << 3;
  assign GEN_3681 = {{1'd0}, T_11934};
  assign T_11974 = GEN_3681 | T_11970;
  assign GEN_3682 = {{4'd0}, pending_36};
  assign T_12010 = GEN_3682 << 4;
  assign GEN_3683 = {{1'd0}, T_11974};
  assign T_12014 = GEN_3683 | T_12010;
  assign GEN_3684 = {{5'd0}, pending_37};
  assign T_12050 = GEN_3684 << 5;
  assign GEN_3685 = {{1'd0}, T_12014};
  assign T_12054 = GEN_3685 | T_12050;
  assign GEN_3686 = {{6'd0}, pending_38};
  assign T_12090 = GEN_3686 << 6;
  assign GEN_3687 = {{1'd0}, T_12054};
  assign T_12094 = GEN_3687 | T_12090;
  assign GEN_3688 = {{7'd0}, pending_39};
  assign T_12130 = GEN_3688 << 7;
  assign GEN_3689 = {{1'd0}, T_12094};
  assign T_12134 = GEN_3689 | T_12130;
  assign GEN_3690 = {{8'd0}, pending_40};
  assign T_12170 = GEN_3690 << 8;
  assign GEN_3691 = {{1'd0}, T_12134};
  assign T_12174 = GEN_3691 | T_12170;
  assign GEN_3692 = {{9'd0}, pending_41};
  assign T_12210 = GEN_3692 << 9;
  assign GEN_3693 = {{1'd0}, T_12174};
  assign T_12214 = GEN_3693 | T_12210;
  assign GEN_3694 = {{10'd0}, pending_42};
  assign T_12250 = GEN_3694 << 10;
  assign GEN_3695 = {{1'd0}, T_12214};
  assign T_12254 = GEN_3695 | T_12250;
  assign GEN_3696 = {{11'd0}, pending_43};
  assign T_12290 = GEN_3696 << 11;
  assign GEN_3697 = {{1'd0}, T_12254};
  assign T_12294 = GEN_3697 | T_12290;
  assign GEN_3698 = {{12'd0}, pending_44};
  assign T_12330 = GEN_3698 << 12;
  assign GEN_3699 = {{1'd0}, T_12294};
  assign T_12334 = GEN_3699 | T_12330;
  assign GEN_3700 = {{13'd0}, pending_45};
  assign T_12370 = GEN_3700 << 13;
  assign GEN_3701 = {{1'd0}, T_12334};
  assign T_12374 = GEN_3701 | T_12370;
  assign GEN_3702 = {{14'd0}, pending_46};
  assign T_12410 = GEN_3702 << 14;
  assign GEN_3703 = {{1'd0}, T_12374};
  assign T_12414 = GEN_3703 | T_12410;
  assign GEN_3704 = {{15'd0}, pending_47};
  assign T_12450 = GEN_3704 << 15;
  assign GEN_3705 = {{1'd0}, T_12414};
  assign T_12454 = GEN_3705 | T_12450;
  assign GEN_3706 = {{16'd0}, pending_48};
  assign T_12490 = GEN_3706 << 16;
  assign GEN_3707 = {{1'd0}, T_12454};
  assign T_12494 = GEN_3707 | T_12490;
  assign GEN_3708 = {{17'd0}, pending_49};
  assign T_12530 = GEN_3708 << 17;
  assign GEN_3709 = {{1'd0}, T_12494};
  assign T_12534 = GEN_3709 | T_12530;
  assign GEN_3710 = {{18'd0}, pending_50};
  assign T_12570 = GEN_3710 << 18;
  assign GEN_3711 = {{1'd0}, T_12534};
  assign T_12574 = GEN_3711 | T_12570;
  assign GEN_3712 = {{19'd0}, pending_51};
  assign T_12610 = GEN_3712 << 19;
  assign GEN_3713 = {{1'd0}, T_12574};
  assign T_12614 = GEN_3713 | T_12610;
  assign T_12634 = T_4344_141 & T_8238;
  assign GEN_406 = T_12634 ? T_3205_bits_data : {{29'd0}, priority_18};
  assign T_12653 = {{29'd0}, priority_18};
  assign T_12674 = T_4344_142 & T_8238;
  assign GEN_407 = T_12674 ? T_3205_bits_data : {{29'd0}, priority_50};
  assign T_12693 = {{29'd0}, priority_50};
  assign T_12714 = T_4344_143 & T_8238;
  assign GEN_408 = T_12714 ? T_3205_bits_data : {{29'd0}, priority_16};
  assign T_12733 = {{29'd0}, priority_16};
  assign T_12754 = T_4344_144 & T_8238;
  assign GEN_409 = T_12754 ? T_3205_bits_data : {{29'd0}, priority_31};
  assign T_12773 = {{29'd0}, priority_31};
  assign T_12794 = T_4344_145 & T_8238;
  assign GEN_410 = T_12794 ? T_3205_bits_data : {{29'd0}, priority_11};
  assign T_12813 = {{29'd0}, priority_11};
  assign T_12834 = T_4344_146 & T_8238;
  assign GEN_411 = T_12834 ? T_3205_bits_data : {{29'd0}, priority_43};
  assign T_12853 = {{29'd0}, priority_43};
  assign T_12874 = T_4344_147 & T_8238;
  assign GEN_412 = T_12874 ? T_3205_bits_data : {{29'd0}, priority_40};
  assign T_12893 = {{29'd0}, priority_40};
  assign T_12914 = T_4344_148 & T_8238;
  assign GEN_413 = T_12914 ? T_3205_bits_data : {{29'd0}, priority_26};
  assign T_12933 = {{29'd0}, priority_26};
  assign T_12954 = T_4344_149 & T_8238;
  assign GEN_414 = T_12954 ? T_3205_bits_data : {{29'd0}, priority_23};
  assign T_12973 = {{29'd0}, priority_23};
  assign T_12994 = T_4344_150 & T_8238;
  assign GEN_415 = T_12994 ? T_3205_bits_data : {{29'd0}, priority_8};
  assign T_13013 = {{29'd0}, priority_8};
  assign T_13034 = T_4344_151 & T_8238;
  assign GEN_416 = T_13034 ? T_3205_bits_data : {{29'd0}, priority_36};
  assign T_13053 = {{29'd0}, priority_36};
  assign T_13074 = T_4344_152 & T_8238;
  assign GEN_417 = T_13074 ? T_3205_bits_data : {{29'd0}, priority_30};
  assign T_13093 = {{29'd0}, priority_30};
  assign T_13114 = T_4344_153 & T_8238;
  assign GEN_418 = T_13114 ? T_3205_bits_data : {{29'd0}, priority_51};
  assign T_13133 = {{29'd0}, priority_51};
  assign T_13154 = T_4344_154 & T_8238;
  assign GEN_419 = T_13154 ? T_3205_bits_data : {{29'd0}, priority_19};
  assign T_13173 = {{29'd0}, priority_19};
  assign T_13194 = T_4344_155 & T_8238;
  assign GEN_420 = T_13194 ? T_3205_bits_data : {{29'd0}, priority_4};
  assign T_13213 = {{29'd0}, priority_4};
  assign T_13234 = T_4344_156 & T_8238;
  assign GEN_421 = T_13234 ? T_3205_bits_data : {{29'd0}, priority_47};
  assign T_13253 = {{29'd0}, priority_47};
  assign T_13274 = T_4344_157 & T_8238;
  assign GEN_422 = T_13274 ? T_3205_bits_data : {{29'd0}, priority_15};
  assign T_13293 = {{29'd0}, priority_15};
  assign T_13541 = T_4319_31 & T_4319_30;
  assign T_13542 = T_13541 & T_4319_29;
  assign T_13543 = T_13542 & T_4319_28;
  assign T_13544 = T_13543 & T_4319_27;
  assign T_13545 = T_13544 & T_4319_26;
  assign T_13546 = T_13545 & T_4319_25;
  assign T_13547 = T_13546 & T_4319_24;
  assign T_13548 = T_13547 & T_4319_23;
  assign T_13549 = T_13548 & T_4319_22;
  assign T_13550 = T_13549 & T_4319_21;
  assign T_13551 = T_13550 & T_4319_20;
  assign T_13552 = T_13551 & T_4319_19;
  assign T_13553 = T_13552 & T_4319_18;
  assign T_13554 = T_13553 & T_4319_17;
  assign T_13555 = T_13554 & T_4319_16;
  assign T_13556 = T_13555 & T_4319_15;
  assign T_13557 = T_13556 & T_4319_14;
  assign T_13558 = T_13557 & T_4319_13;
  assign T_13559 = T_13558 & T_4319_12;
  assign T_13560 = T_13559 & T_4319_11;
  assign T_13561 = T_13560 & T_4319_10;
  assign T_13562 = T_13561 & T_4319_9;
  assign T_13563 = T_13562 & T_4319_8;
  assign T_13564 = T_13563 & T_4319_7;
  assign T_13565 = T_13564 & T_4319_6;
  assign T_13566 = T_13565 & T_4319_5;
  assign T_13567 = T_13566 & T_4319_4;
  assign T_13568 = T_13567 & T_4319_3;
  assign T_13569 = T_13568 & T_4319_2;
  assign T_13570 = T_13569 & T_4319_1;
  assign T_13571 = T_13570 & T_4319_0;
  assign T_13576 = T_4319_140 & T_4319_139;
  assign T_13577 = T_13576 & T_4319_138;
  assign T_13578 = T_13577 & T_4319_137;
  assign T_13579 = T_13578 & T_4319_136;
  assign T_13580 = T_13579 & T_4319_135;
  assign T_13581 = T_13580 & T_4319_134;
  assign T_13582 = T_13581 & T_4319_133;
  assign T_13583 = T_13582 & T_4319_132;
  assign T_13584 = T_13583 & T_4319_131;
  assign T_13585 = T_13584 & T_4319_130;
  assign T_13586 = T_13585 & T_4319_129;
  assign T_13587 = T_13586 & T_4319_128;
  assign T_13588 = T_13587 & T_4319_127;
  assign T_13589 = T_13588 & T_4319_126;
  assign T_13590 = T_13589 & T_4319_125;
  assign T_13591 = T_13590 & T_4319_124;
  assign T_13592 = T_13591 & T_4319_123;
  assign T_13593 = T_13592 & T_4319_122;
  assign T_13594 = T_13593 & T_4319_121;
  assign T_13785 = T_4319_110 & T_4319_109;
  assign T_13786 = T_13785 & T_4319_108;
  assign T_13787 = T_13786 & T_4319_107;
  assign T_13788 = T_13787 & T_4319_106;
  assign T_13789 = T_13788 & T_4319_105;
  assign T_13790 = T_13789 & T_4319_104;
  assign T_13791 = T_13790 & T_4319_103;
  assign T_13792 = T_13791 & T_4319_102;
  assign T_13793 = T_13792 & T_4319_101;
  assign T_13794 = T_13793 & T_4319_100;
  assign T_13795 = T_13794 & T_4319_99;
  assign T_13796 = T_13795 & T_4319_98;
  assign T_13797 = T_13796 & T_4319_97;
  assign T_13798 = T_13797 & T_4319_96;
  assign T_13799 = T_13798 & T_4319_95;
  assign T_13800 = T_13799 & T_4319_94;
  assign T_13801 = T_13800 & T_4319_93;
  assign T_13802 = T_13801 & T_4319_92;
  assign T_13803 = T_13802 & T_4319_91;
  assign T_13804 = T_13803 & T_4319_90;
  assign T_13805 = T_13804 & T_4319_89;
  assign T_13806 = T_13805 & T_4319_88;
  assign T_13807 = T_13806 & T_4319_87;
  assign T_13808 = T_13807 & T_4319_86;
  assign T_13809 = T_13808 & T_4319_85;
  assign T_13810 = T_13809 & T_4319_84;
  assign T_13811 = T_13810 & T_4319_83;
  assign T_13812 = T_13811 & T_4319_82;
  assign T_13813 = T_13812 & T_4319_81;
  assign T_13814 = T_13813 & T_4319_80;
  assign T_13815 = T_13814 & T_4319_79;
  assign T_13820 = T_4319_60 & T_4319_59;
  assign T_13821 = T_13820 & T_4319_58;
  assign T_13822 = T_13821 & T_4319_57;
  assign T_13823 = T_13822 & T_4319_56;
  assign T_13824 = T_13823 & T_4319_55;
  assign T_13825 = T_13824 & T_4319_54;
  assign T_13826 = T_13825 & T_4319_53;
  assign T_13827 = T_13826 & T_4319_52;
  assign T_13828 = T_13827 & T_4319_51;
  assign T_13829 = T_13828 & T_4319_50;
  assign T_13830 = T_13829 & T_4319_49;
  assign T_13831 = T_13830 & T_4319_48;
  assign T_13832 = T_13831 & T_4319_47;
  assign T_13833 = T_13832 & T_4319_46;
  assign T_13834 = T_13833 & T_4319_45;
  assign T_13835 = T_13834 & T_4319_44;
  assign T_13836 = T_13835 & T_4319_43;
  assign T_13837 = T_13836 & T_4319_42;
  assign T_13838 = T_13837 & T_4319_41;
  assign T_15504_0 = T_4319_32;
  assign T_15504_1 = T_4319_64;
  assign T_15504_2 = T_4319_73;
  assign T_15504_3 = T_4319_118;
  assign T_15504_4 = T_4319_155;
  assign T_15504_5 = T_4319_33;
  assign T_15504_6 = T_4319_65;
  assign T_15504_7 = T_4319_116;
  assign T_15504_8 = T_4319_150;
  assign T_15504_9 = T_4319_70;
  assign T_15504_10 = T_4319_34;
  assign T_15504_11 = T_4319_145;
  assign T_15504_12 = T_4319_114;
  assign T_15504_13 = T_4319_71;
  assign T_15504_14 = T_4319_39;
  assign T_15504_15 = T_4319_157;
  assign T_15504_16 = T_4319_143;
  assign T_15504_17 = T_4319_77;
  assign T_15504_18 = T_4319_141;
  assign T_15504_19 = T_4319_154;
  assign T_15504_20 = T_4319_40;
  assign T_15504_21 = T_4319_68;
  assign T_15504_22 = T_4319_111;
  assign T_15504_23 = T_4319_149;
  assign T_15504_24 = T_4319_36;
  assign T_15504_25 = T_4319_38;
  assign T_15504_26 = T_4319_148;
  assign T_15504_27 = T_4319_113;
  assign T_15504_28 = T_4319_66;
  assign T_15504_29 = T_4319_62;
  assign T_15504_30 = T_4319_152;
  assign T_15504_31 = T_4319_144;
  assign T_15504_32 = T_4319_74;
  assign T_15504_33 = T_4319_69;
  assign T_15504_34 = T_4319_75;
  assign T_15504_35 = T_4319_119;
  assign T_15504_36 = T_4319_151;
  assign T_15504_37 = T_4319_37;
  assign T_15504_38 = T_4319_67;
  assign T_15504_39 = T_4319_117;
  assign T_15504_40 = T_4319_147;
  assign T_15504_41 = T_4319_72;
  assign T_15504_42 = T_4319_35;
  assign T_15504_43 = T_4319_146;
  assign T_15504_44 = T_4319_112;
  assign T_15504_45 = T_4319_76;
  assign T_15504_46 = T_4319_61;
  assign T_15504_47 = T_4319_156;
  assign T_15504_48 = T_4319_120;
  assign T_15504_49 = T_4319_115;
  assign T_15504_50 = T_4319_142;
  assign T_15504_51 = T_4319_153;
  assign T_15504_52 = 1'h1;
  assign T_15504_53 = 1'h1;
  assign T_15504_54 = 1'h1;
  assign T_15504_55 = 1'h1;
  assign T_15504_56 = 1'h1;
  assign T_15504_57 = 1'h1;
  assign T_15504_58 = 1'h1;
  assign T_15504_59 = 1'h1;
  assign T_15504_60 = 1'h1;
  assign T_15504_61 = 1'h1;
  assign T_15504_62 = 1'h1;
  assign T_15504_63 = 1'h1;
  assign T_15504_64 = T_13571;
  assign T_15504_65 = T_13594;
  assign T_15504_66 = 1'h1;
  assign T_15504_67 = 1'h1;
  assign T_15504_68 = 1'h1;
  assign T_15504_69 = 1'h1;
  assign T_15504_70 = 1'h1;
  assign T_15504_71 = 1'h1;
  assign T_15504_72 = 1'h1;
  assign T_15504_73 = 1'h1;
  assign T_15504_74 = 1'h1;
  assign T_15504_75 = 1'h1;
  assign T_15504_76 = 1'h1;
  assign T_15504_77 = 1'h1;
  assign T_15504_78 = 1'h1;
  assign T_15504_79 = 1'h1;
  assign T_15504_80 = 1'h1;
  assign T_15504_81 = 1'h1;
  assign T_15504_82 = 1'h1;
  assign T_15504_83 = 1'h1;
  assign T_15504_84 = 1'h1;
  assign T_15504_85 = 1'h1;
  assign T_15504_86 = 1'h1;
  assign T_15504_87 = 1'h1;
  assign T_15504_88 = 1'h1;
  assign T_15504_89 = 1'h1;
  assign T_15504_90 = 1'h1;
  assign T_15504_91 = 1'h1;
  assign T_15504_92 = 1'h1;
  assign T_15504_93 = 1'h1;
  assign T_15504_94 = 1'h1;
  assign T_15504_95 = 1'h1;
  assign T_15504_96 = 1'h1;
  assign T_15504_97 = 1'h1;
  assign T_15504_98 = 1'h1;
  assign T_15504_99 = 1'h1;
  assign T_15504_100 = 1'h1;
  assign T_15504_101 = 1'h1;
  assign T_15504_102 = 1'h1;
  assign T_15504_103 = 1'h1;
  assign T_15504_104 = 1'h1;
  assign T_15504_105 = 1'h1;
  assign T_15504_106 = 1'h1;
  assign T_15504_107 = 1'h1;
  assign T_15504_108 = 1'h1;
  assign T_15504_109 = 1'h1;
  assign T_15504_110 = 1'h1;
  assign T_15504_111 = 1'h1;
  assign T_15504_112 = 1'h1;
  assign T_15504_113 = 1'h1;
  assign T_15504_114 = 1'h1;
  assign T_15504_115 = 1'h1;
  assign T_15504_116 = 1'h1;
  assign T_15504_117 = 1'h1;
  assign T_15504_118 = 1'h1;
  assign T_15504_119 = 1'h1;
  assign T_15504_120 = 1'h1;
  assign T_15504_121 = 1'h1;
  assign T_15504_122 = 1'h1;
  assign T_15504_123 = 1'h1;
  assign T_15504_124 = 1'h1;
  assign T_15504_125 = 1'h1;
  assign T_15504_126 = 1'h1;
  assign T_15504_127 = 1'h1;
  assign T_15504_128 = T_13815;
  assign T_15504_129 = T_13838;
  assign T_15504_130 = 1'h1;
  assign T_15504_131 = 1'h1;
  assign T_15504_132 = 1'h1;
  assign T_15504_133 = 1'h1;
  assign T_15504_134 = 1'h1;
  assign T_15504_135 = 1'h1;
  assign T_15504_136 = 1'h1;
  assign T_15504_137 = 1'h1;
  assign T_15504_138 = 1'h1;
  assign T_15504_139 = 1'h1;
  assign T_15504_140 = 1'h1;
  assign T_15504_141 = 1'h1;
  assign T_15504_142 = 1'h1;
  assign T_15504_143 = 1'h1;
  assign T_15504_144 = 1'h1;
  assign T_15504_145 = 1'h1;
  assign T_15504_146 = 1'h1;
  assign T_15504_147 = 1'h1;
  assign T_15504_148 = 1'h1;
  assign T_15504_149 = 1'h1;
  assign T_15504_150 = 1'h1;
  assign T_15504_151 = 1'h1;
  assign T_15504_152 = 1'h1;
  assign T_15504_153 = 1'h1;
  assign T_15504_154 = 1'h1;
  assign T_15504_155 = 1'h1;
  assign T_15504_156 = 1'h1;
  assign T_15504_157 = 1'h1;
  assign T_15504_158 = 1'h1;
  assign T_15504_159 = 1'h1;
  assign T_15504_160 = 1'h1;
  assign T_15504_161 = 1'h1;
  assign T_15504_162 = 1'h1;
  assign T_15504_163 = 1'h1;
  assign T_15504_164 = 1'h1;
  assign T_15504_165 = 1'h1;
  assign T_15504_166 = 1'h1;
  assign T_15504_167 = 1'h1;
  assign T_15504_168 = 1'h1;
  assign T_15504_169 = 1'h1;
  assign T_15504_170 = 1'h1;
  assign T_15504_171 = 1'h1;
  assign T_15504_172 = 1'h1;
  assign T_15504_173 = 1'h1;
  assign T_15504_174 = 1'h1;
  assign T_15504_175 = 1'h1;
  assign T_15504_176 = 1'h1;
  assign T_15504_177 = 1'h1;
  assign T_15504_178 = 1'h1;
  assign T_15504_179 = 1'h1;
  assign T_15504_180 = 1'h1;
  assign T_15504_181 = 1'h1;
  assign T_15504_182 = 1'h1;
  assign T_15504_183 = 1'h1;
  assign T_15504_184 = 1'h1;
  assign T_15504_185 = 1'h1;
  assign T_15504_186 = 1'h1;
  assign T_15504_187 = 1'h1;
  assign T_15504_188 = 1'h1;
  assign T_15504_189 = 1'h1;
  assign T_15504_190 = 1'h1;
  assign T_15504_191 = 1'h1;
  assign T_15504_192 = 1'h1;
  assign T_15504_193 = 1'h1;
  assign T_15504_194 = 1'h1;
  assign T_15504_195 = 1'h1;
  assign T_15504_196 = 1'h1;
  assign T_15504_197 = 1'h1;
  assign T_15504_198 = 1'h1;
  assign T_15504_199 = 1'h1;
  assign T_15504_200 = 1'h1;
  assign T_15504_201 = 1'h1;
  assign T_15504_202 = 1'h1;
  assign T_15504_203 = 1'h1;
  assign T_15504_204 = 1'h1;
  assign T_15504_205 = 1'h1;
  assign T_15504_206 = 1'h1;
  assign T_15504_207 = 1'h1;
  assign T_15504_208 = 1'h1;
  assign T_15504_209 = 1'h1;
  assign T_15504_210 = 1'h1;
  assign T_15504_211 = 1'h1;
  assign T_15504_212 = 1'h1;
  assign T_15504_213 = 1'h1;
  assign T_15504_214 = 1'h1;
  assign T_15504_215 = 1'h1;
  assign T_15504_216 = 1'h1;
  assign T_15504_217 = 1'h1;
  assign T_15504_218 = 1'h1;
  assign T_15504_219 = 1'h1;
  assign T_15504_220 = 1'h1;
  assign T_15504_221 = 1'h1;
  assign T_15504_222 = 1'h1;
  assign T_15504_223 = 1'h1;
  assign T_15504_224 = 1'h1;
  assign T_15504_225 = 1'h1;
  assign T_15504_226 = 1'h1;
  assign T_15504_227 = 1'h1;
  assign T_15504_228 = 1'h1;
  assign T_15504_229 = 1'h1;
  assign T_15504_230 = 1'h1;
  assign T_15504_231 = 1'h1;
  assign T_15504_232 = 1'h1;
  assign T_15504_233 = 1'h1;
  assign T_15504_234 = 1'h1;
  assign T_15504_235 = 1'h1;
  assign T_15504_236 = 1'h1;
  assign T_15504_237 = 1'h1;
  assign T_15504_238 = 1'h1;
  assign T_15504_239 = 1'h1;
  assign T_15504_240 = 1'h1;
  assign T_15504_241 = 1'h1;
  assign T_15504_242 = 1'h1;
  assign T_15504_243 = 1'h1;
  assign T_15504_244 = 1'h1;
  assign T_15504_245 = 1'h1;
  assign T_15504_246 = 1'h1;
  assign T_15504_247 = 1'h1;
  assign T_15504_248 = 1'h1;
  assign T_15504_249 = 1'h1;
  assign T_15504_250 = 1'h1;
  assign T_15504_251 = 1'h1;
  assign T_15504_252 = 1'h1;
  assign T_15504_253 = 1'h1;
  assign T_15504_254 = 1'h1;
  assign T_15504_255 = 1'h1;
  assign T_15504_256 = T_4319_78;
  assign T_15504_257 = T_4319_63;
  assign T_15504_258 = 1'h1;
  assign T_15504_259 = 1'h1;
  assign T_15504_260 = 1'h1;
  assign T_15504_261 = 1'h1;
  assign T_15504_262 = 1'h1;
  assign T_15504_263 = 1'h1;
  assign T_15504_264 = 1'h1;
  assign T_15504_265 = 1'h1;
  assign T_15504_266 = 1'h1;
  assign T_15504_267 = 1'h1;
  assign T_15504_268 = 1'h1;
  assign T_15504_269 = 1'h1;
  assign T_15504_270 = 1'h1;
  assign T_15504_271 = 1'h1;
  assign T_15504_272 = 1'h1;
  assign T_15504_273 = 1'h1;
  assign T_15504_274 = 1'h1;
  assign T_15504_275 = 1'h1;
  assign T_15504_276 = 1'h1;
  assign T_15504_277 = 1'h1;
  assign T_15504_278 = 1'h1;
  assign T_15504_279 = 1'h1;
  assign T_15504_280 = 1'h1;
  assign T_15504_281 = 1'h1;
  assign T_15504_282 = 1'h1;
  assign T_15504_283 = 1'h1;
  assign T_15504_284 = 1'h1;
  assign T_15504_285 = 1'h1;
  assign T_15504_286 = 1'h1;
  assign T_15504_287 = 1'h1;
  assign T_15504_288 = 1'h1;
  assign T_15504_289 = 1'h1;
  assign T_15504_290 = 1'h1;
  assign T_15504_291 = 1'h1;
  assign T_15504_292 = 1'h1;
  assign T_15504_293 = 1'h1;
  assign T_15504_294 = 1'h1;
  assign T_15504_295 = 1'h1;
  assign T_15504_296 = 1'h1;
  assign T_15504_297 = 1'h1;
  assign T_15504_298 = 1'h1;
  assign T_15504_299 = 1'h1;
  assign T_15504_300 = 1'h1;
  assign T_15504_301 = 1'h1;
  assign T_15504_302 = 1'h1;
  assign T_15504_303 = 1'h1;
  assign T_15504_304 = 1'h1;
  assign T_15504_305 = 1'h1;
  assign T_15504_306 = 1'h1;
  assign T_15504_307 = 1'h1;
  assign T_15504_308 = 1'h1;
  assign T_15504_309 = 1'h1;
  assign T_15504_310 = 1'h1;
  assign T_15504_311 = 1'h1;
  assign T_15504_312 = 1'h1;
  assign T_15504_313 = 1'h1;
  assign T_15504_314 = 1'h1;
  assign T_15504_315 = 1'h1;
  assign T_15504_316 = 1'h1;
  assign T_15504_317 = 1'h1;
  assign T_15504_318 = 1'h1;
  assign T_15504_319 = 1'h1;
  assign T_15504_320 = 1'h1;
  assign T_15504_321 = 1'h1;
  assign T_15504_322 = 1'h1;
  assign T_15504_323 = 1'h1;
  assign T_15504_324 = 1'h1;
  assign T_15504_325 = 1'h1;
  assign T_15504_326 = 1'h1;
  assign T_15504_327 = 1'h1;
  assign T_15504_328 = 1'h1;
  assign T_15504_329 = 1'h1;
  assign T_15504_330 = 1'h1;
  assign T_15504_331 = 1'h1;
  assign T_15504_332 = 1'h1;
  assign T_15504_333 = 1'h1;
  assign T_15504_334 = 1'h1;
  assign T_15504_335 = 1'h1;
  assign T_15504_336 = 1'h1;
  assign T_15504_337 = 1'h1;
  assign T_15504_338 = 1'h1;
  assign T_15504_339 = 1'h1;
  assign T_15504_340 = 1'h1;
  assign T_15504_341 = 1'h1;
  assign T_15504_342 = 1'h1;
  assign T_15504_343 = 1'h1;
  assign T_15504_344 = 1'h1;
  assign T_15504_345 = 1'h1;
  assign T_15504_346 = 1'h1;
  assign T_15504_347 = 1'h1;
  assign T_15504_348 = 1'h1;
  assign T_15504_349 = 1'h1;
  assign T_15504_350 = 1'h1;
  assign T_15504_351 = 1'h1;
  assign T_15504_352 = 1'h1;
  assign T_15504_353 = 1'h1;
  assign T_15504_354 = 1'h1;
  assign T_15504_355 = 1'h1;
  assign T_15504_356 = 1'h1;
  assign T_15504_357 = 1'h1;
  assign T_15504_358 = 1'h1;
  assign T_15504_359 = 1'h1;
  assign T_15504_360 = 1'h1;
  assign T_15504_361 = 1'h1;
  assign T_15504_362 = 1'h1;
  assign T_15504_363 = 1'h1;
  assign T_15504_364 = 1'h1;
  assign T_15504_365 = 1'h1;
  assign T_15504_366 = 1'h1;
  assign T_15504_367 = 1'h1;
  assign T_15504_368 = 1'h1;
  assign T_15504_369 = 1'h1;
  assign T_15504_370 = 1'h1;
  assign T_15504_371 = 1'h1;
  assign T_15504_372 = 1'h1;
  assign T_15504_373 = 1'h1;
  assign T_15504_374 = 1'h1;
  assign T_15504_375 = 1'h1;
  assign T_15504_376 = 1'h1;
  assign T_15504_377 = 1'h1;
  assign T_15504_378 = 1'h1;
  assign T_15504_379 = 1'h1;
  assign T_15504_380 = 1'h1;
  assign T_15504_381 = 1'h1;
  assign T_15504_382 = 1'h1;
  assign T_15504_383 = 1'h1;
  assign T_15504_384 = 1'h1;
  assign T_15504_385 = 1'h1;
  assign T_15504_386 = 1'h1;
  assign T_15504_387 = 1'h1;
  assign T_15504_388 = 1'h1;
  assign T_15504_389 = 1'h1;
  assign T_15504_390 = 1'h1;
  assign T_15504_391 = 1'h1;
  assign T_15504_392 = 1'h1;
  assign T_15504_393 = 1'h1;
  assign T_15504_394 = 1'h1;
  assign T_15504_395 = 1'h1;
  assign T_15504_396 = 1'h1;
  assign T_15504_397 = 1'h1;
  assign T_15504_398 = 1'h1;
  assign T_15504_399 = 1'h1;
  assign T_15504_400 = 1'h1;
  assign T_15504_401 = 1'h1;
  assign T_15504_402 = 1'h1;
  assign T_15504_403 = 1'h1;
  assign T_15504_404 = 1'h1;
  assign T_15504_405 = 1'h1;
  assign T_15504_406 = 1'h1;
  assign T_15504_407 = 1'h1;
  assign T_15504_408 = 1'h1;
  assign T_15504_409 = 1'h1;
  assign T_15504_410 = 1'h1;
  assign T_15504_411 = 1'h1;
  assign T_15504_412 = 1'h1;
  assign T_15504_413 = 1'h1;
  assign T_15504_414 = 1'h1;
  assign T_15504_415 = 1'h1;
  assign T_15504_416 = 1'h1;
  assign T_15504_417 = 1'h1;
  assign T_15504_418 = 1'h1;
  assign T_15504_419 = 1'h1;
  assign T_15504_420 = 1'h1;
  assign T_15504_421 = 1'h1;
  assign T_15504_422 = 1'h1;
  assign T_15504_423 = 1'h1;
  assign T_15504_424 = 1'h1;
  assign T_15504_425 = 1'h1;
  assign T_15504_426 = 1'h1;
  assign T_15504_427 = 1'h1;
  assign T_15504_428 = 1'h1;
  assign T_15504_429 = 1'h1;
  assign T_15504_430 = 1'h1;
  assign T_15504_431 = 1'h1;
  assign T_15504_432 = 1'h1;
  assign T_15504_433 = 1'h1;
  assign T_15504_434 = 1'h1;
  assign T_15504_435 = 1'h1;
  assign T_15504_436 = 1'h1;
  assign T_15504_437 = 1'h1;
  assign T_15504_438 = 1'h1;
  assign T_15504_439 = 1'h1;
  assign T_15504_440 = 1'h1;
  assign T_15504_441 = 1'h1;
  assign T_15504_442 = 1'h1;
  assign T_15504_443 = 1'h1;
  assign T_15504_444 = 1'h1;
  assign T_15504_445 = 1'h1;
  assign T_15504_446 = 1'h1;
  assign T_15504_447 = 1'h1;
  assign T_15504_448 = 1'h1;
  assign T_15504_449 = 1'h1;
  assign T_15504_450 = 1'h1;
  assign T_15504_451 = 1'h1;
  assign T_15504_452 = 1'h1;
  assign T_15504_453 = 1'h1;
  assign T_15504_454 = 1'h1;
  assign T_15504_455 = 1'h1;
  assign T_15504_456 = 1'h1;
  assign T_15504_457 = 1'h1;
  assign T_15504_458 = 1'h1;
  assign T_15504_459 = 1'h1;
  assign T_15504_460 = 1'h1;
  assign T_15504_461 = 1'h1;
  assign T_15504_462 = 1'h1;
  assign T_15504_463 = 1'h1;
  assign T_15504_464 = 1'h1;
  assign T_15504_465 = 1'h1;
  assign T_15504_466 = 1'h1;
  assign T_15504_467 = 1'h1;
  assign T_15504_468 = 1'h1;
  assign T_15504_469 = 1'h1;
  assign T_15504_470 = 1'h1;
  assign T_15504_471 = 1'h1;
  assign T_15504_472 = 1'h1;
  assign T_15504_473 = 1'h1;
  assign T_15504_474 = 1'h1;
  assign T_15504_475 = 1'h1;
  assign T_15504_476 = 1'h1;
  assign T_15504_477 = 1'h1;
  assign T_15504_478 = 1'h1;
  assign T_15504_479 = 1'h1;
  assign T_15504_480 = 1'h1;
  assign T_15504_481 = 1'h1;
  assign T_15504_482 = 1'h1;
  assign T_15504_483 = 1'h1;
  assign T_15504_484 = 1'h1;
  assign T_15504_485 = 1'h1;
  assign T_15504_486 = 1'h1;
  assign T_15504_487 = 1'h1;
  assign T_15504_488 = 1'h1;
  assign T_15504_489 = 1'h1;
  assign T_15504_490 = 1'h1;
  assign T_15504_491 = 1'h1;
  assign T_15504_492 = 1'h1;
  assign T_15504_493 = 1'h1;
  assign T_15504_494 = 1'h1;
  assign T_15504_495 = 1'h1;
  assign T_15504_496 = 1'h1;
  assign T_15504_497 = 1'h1;
  assign T_15504_498 = 1'h1;
  assign T_15504_499 = 1'h1;
  assign T_15504_500 = 1'h1;
  assign T_15504_501 = 1'h1;
  assign T_15504_502 = 1'h1;
  assign T_15504_503 = 1'h1;
  assign T_15504_504 = 1'h1;
  assign T_15504_505 = 1'h1;
  assign T_15504_506 = 1'h1;
  assign T_15504_507 = 1'h1;
  assign T_15504_508 = 1'h1;
  assign T_15504_509 = 1'h1;
  assign T_15504_510 = 1'h1;
  assign T_15504_511 = 1'h1;
  assign T_16265 = T_4324_31 & T_4324_30;
  assign T_16266 = T_16265 & T_4324_29;
  assign T_16267 = T_16266 & T_4324_28;
  assign T_16268 = T_16267 & T_4324_27;
  assign T_16269 = T_16268 & T_4324_26;
  assign T_16270 = T_16269 & T_4324_25;
  assign T_16271 = T_16270 & T_4324_24;
  assign T_16272 = T_16271 & T_4324_23;
  assign T_16273 = T_16272 & T_4324_22;
  assign T_16274 = T_16273 & T_4324_21;
  assign T_16275 = T_16274 & T_4324_20;
  assign T_16276 = T_16275 & T_4324_19;
  assign T_16277 = T_16276 & T_4324_18;
  assign T_16278 = T_16277 & T_4324_17;
  assign T_16279 = T_16278 & T_4324_16;
  assign T_16280 = T_16279 & T_4324_15;
  assign T_16281 = T_16280 & T_4324_14;
  assign T_16282 = T_16281 & T_4324_13;
  assign T_16283 = T_16282 & T_4324_12;
  assign T_16284 = T_16283 & T_4324_11;
  assign T_16285 = T_16284 & T_4324_10;
  assign T_16286 = T_16285 & T_4324_9;
  assign T_16287 = T_16286 & T_4324_8;
  assign T_16288 = T_16287 & T_4324_7;
  assign T_16289 = T_16288 & T_4324_6;
  assign T_16290 = T_16289 & T_4324_5;
  assign T_16291 = T_16290 & T_4324_4;
  assign T_16292 = T_16291 & T_4324_3;
  assign T_16293 = T_16292 & T_4324_2;
  assign T_16294 = T_16293 & T_4324_1;
  assign T_16295 = T_16294 & T_4324_0;
  assign T_16300 = T_4324_140 & T_4324_139;
  assign T_16301 = T_16300 & T_4324_138;
  assign T_16302 = T_16301 & T_4324_137;
  assign T_16303 = T_16302 & T_4324_136;
  assign T_16304 = T_16303 & T_4324_135;
  assign T_16305 = T_16304 & T_4324_134;
  assign T_16306 = T_16305 & T_4324_133;
  assign T_16307 = T_16306 & T_4324_132;
  assign T_16308 = T_16307 & T_4324_131;
  assign T_16309 = T_16308 & T_4324_130;
  assign T_16310 = T_16309 & T_4324_129;
  assign T_16311 = T_16310 & T_4324_128;
  assign T_16312 = T_16311 & T_4324_127;
  assign T_16313 = T_16312 & T_4324_126;
  assign T_16314 = T_16313 & T_4324_125;
  assign T_16315 = T_16314 & T_4324_124;
  assign T_16316 = T_16315 & T_4324_123;
  assign T_16317 = T_16316 & T_4324_122;
  assign T_16318 = T_16317 & T_4324_121;
  assign T_16509 = T_4324_110 & T_4324_109;
  assign T_16510 = T_16509 & T_4324_108;
  assign T_16511 = T_16510 & T_4324_107;
  assign T_16512 = T_16511 & T_4324_106;
  assign T_16513 = T_16512 & T_4324_105;
  assign T_16514 = T_16513 & T_4324_104;
  assign T_16515 = T_16514 & T_4324_103;
  assign T_16516 = T_16515 & T_4324_102;
  assign T_16517 = T_16516 & T_4324_101;
  assign T_16518 = T_16517 & T_4324_100;
  assign T_16519 = T_16518 & T_4324_99;
  assign T_16520 = T_16519 & T_4324_98;
  assign T_16521 = T_16520 & T_4324_97;
  assign T_16522 = T_16521 & T_4324_96;
  assign T_16523 = T_16522 & T_4324_95;
  assign T_16524 = T_16523 & T_4324_94;
  assign T_16525 = T_16524 & T_4324_93;
  assign T_16526 = T_16525 & T_4324_92;
  assign T_16527 = T_16526 & T_4324_91;
  assign T_16528 = T_16527 & T_4324_90;
  assign T_16529 = T_16528 & T_4324_89;
  assign T_16530 = T_16529 & T_4324_88;
  assign T_16531 = T_16530 & T_4324_87;
  assign T_16532 = T_16531 & T_4324_86;
  assign T_16533 = T_16532 & T_4324_85;
  assign T_16534 = T_16533 & T_4324_84;
  assign T_16535 = T_16534 & T_4324_83;
  assign T_16536 = T_16535 & T_4324_82;
  assign T_16537 = T_16536 & T_4324_81;
  assign T_16538 = T_16537 & T_4324_80;
  assign T_16539 = T_16538 & T_4324_79;
  assign T_16544 = T_4324_60 & T_4324_59;
  assign T_16545 = T_16544 & T_4324_58;
  assign T_16546 = T_16545 & T_4324_57;
  assign T_16547 = T_16546 & T_4324_56;
  assign T_16548 = T_16547 & T_4324_55;
  assign T_16549 = T_16548 & T_4324_54;
  assign T_16550 = T_16549 & T_4324_53;
  assign T_16551 = T_16550 & T_4324_52;
  assign T_16552 = T_16551 & T_4324_51;
  assign T_16553 = T_16552 & T_4324_50;
  assign T_16554 = T_16553 & T_4324_49;
  assign T_16555 = T_16554 & T_4324_48;
  assign T_16556 = T_16555 & T_4324_47;
  assign T_16557 = T_16556 & T_4324_46;
  assign T_16558 = T_16557 & T_4324_45;
  assign T_16559 = T_16558 & T_4324_44;
  assign T_16560 = T_16559 & T_4324_43;
  assign T_16561 = T_16560 & T_4324_42;
  assign T_16562 = T_16561 & T_4324_41;
  assign T_18228_0 = T_4324_32;
  assign T_18228_1 = T_4324_64;
  assign T_18228_2 = T_4324_73;
  assign T_18228_3 = T_4324_118;
  assign T_18228_4 = T_4324_155;
  assign T_18228_5 = T_4324_33;
  assign T_18228_6 = T_4324_65;
  assign T_18228_7 = T_4324_116;
  assign T_18228_8 = T_4324_150;
  assign T_18228_9 = T_4324_70;
  assign T_18228_10 = T_4324_34;
  assign T_18228_11 = T_4324_145;
  assign T_18228_12 = T_4324_114;
  assign T_18228_13 = T_4324_71;
  assign T_18228_14 = T_4324_39;
  assign T_18228_15 = T_4324_157;
  assign T_18228_16 = T_4324_143;
  assign T_18228_17 = T_4324_77;
  assign T_18228_18 = T_4324_141;
  assign T_18228_19 = T_4324_154;
  assign T_18228_20 = T_4324_40;
  assign T_18228_21 = T_4324_68;
  assign T_18228_22 = T_4324_111;
  assign T_18228_23 = T_4324_149;
  assign T_18228_24 = T_4324_36;
  assign T_18228_25 = T_4324_38;
  assign T_18228_26 = T_4324_148;
  assign T_18228_27 = T_4324_113;
  assign T_18228_28 = T_4324_66;
  assign T_18228_29 = T_4324_62;
  assign T_18228_30 = T_4324_152;
  assign T_18228_31 = T_4324_144;
  assign T_18228_32 = T_4324_74;
  assign T_18228_33 = T_4324_69;
  assign T_18228_34 = T_4324_75;
  assign T_18228_35 = T_4324_119;
  assign T_18228_36 = T_4324_151;
  assign T_18228_37 = T_4324_37;
  assign T_18228_38 = T_4324_67;
  assign T_18228_39 = T_4324_117;
  assign T_18228_40 = T_4324_147;
  assign T_18228_41 = T_4324_72;
  assign T_18228_42 = T_4324_35;
  assign T_18228_43 = T_4324_146;
  assign T_18228_44 = T_4324_112;
  assign T_18228_45 = T_4324_76;
  assign T_18228_46 = T_4324_61;
  assign T_18228_47 = T_4324_156;
  assign T_18228_48 = T_4324_120;
  assign T_18228_49 = T_4324_115;
  assign T_18228_50 = T_4324_142;
  assign T_18228_51 = T_4324_153;
  assign T_18228_52 = 1'h1;
  assign T_18228_53 = 1'h1;
  assign T_18228_54 = 1'h1;
  assign T_18228_55 = 1'h1;
  assign T_18228_56 = 1'h1;
  assign T_18228_57 = 1'h1;
  assign T_18228_58 = 1'h1;
  assign T_18228_59 = 1'h1;
  assign T_18228_60 = 1'h1;
  assign T_18228_61 = 1'h1;
  assign T_18228_62 = 1'h1;
  assign T_18228_63 = 1'h1;
  assign T_18228_64 = T_16295;
  assign T_18228_65 = T_16318;
  assign T_18228_66 = 1'h1;
  assign T_18228_67 = 1'h1;
  assign T_18228_68 = 1'h1;
  assign T_18228_69 = 1'h1;
  assign T_18228_70 = 1'h1;
  assign T_18228_71 = 1'h1;
  assign T_18228_72 = 1'h1;
  assign T_18228_73 = 1'h1;
  assign T_18228_74 = 1'h1;
  assign T_18228_75 = 1'h1;
  assign T_18228_76 = 1'h1;
  assign T_18228_77 = 1'h1;
  assign T_18228_78 = 1'h1;
  assign T_18228_79 = 1'h1;
  assign T_18228_80 = 1'h1;
  assign T_18228_81 = 1'h1;
  assign T_18228_82 = 1'h1;
  assign T_18228_83 = 1'h1;
  assign T_18228_84 = 1'h1;
  assign T_18228_85 = 1'h1;
  assign T_18228_86 = 1'h1;
  assign T_18228_87 = 1'h1;
  assign T_18228_88 = 1'h1;
  assign T_18228_89 = 1'h1;
  assign T_18228_90 = 1'h1;
  assign T_18228_91 = 1'h1;
  assign T_18228_92 = 1'h1;
  assign T_18228_93 = 1'h1;
  assign T_18228_94 = 1'h1;
  assign T_18228_95 = 1'h1;
  assign T_18228_96 = 1'h1;
  assign T_18228_97 = 1'h1;
  assign T_18228_98 = 1'h1;
  assign T_18228_99 = 1'h1;
  assign T_18228_100 = 1'h1;
  assign T_18228_101 = 1'h1;
  assign T_18228_102 = 1'h1;
  assign T_18228_103 = 1'h1;
  assign T_18228_104 = 1'h1;
  assign T_18228_105 = 1'h1;
  assign T_18228_106 = 1'h1;
  assign T_18228_107 = 1'h1;
  assign T_18228_108 = 1'h1;
  assign T_18228_109 = 1'h1;
  assign T_18228_110 = 1'h1;
  assign T_18228_111 = 1'h1;
  assign T_18228_112 = 1'h1;
  assign T_18228_113 = 1'h1;
  assign T_18228_114 = 1'h1;
  assign T_18228_115 = 1'h1;
  assign T_18228_116 = 1'h1;
  assign T_18228_117 = 1'h1;
  assign T_18228_118 = 1'h1;
  assign T_18228_119 = 1'h1;
  assign T_18228_120 = 1'h1;
  assign T_18228_121 = 1'h1;
  assign T_18228_122 = 1'h1;
  assign T_18228_123 = 1'h1;
  assign T_18228_124 = 1'h1;
  assign T_18228_125 = 1'h1;
  assign T_18228_126 = 1'h1;
  assign T_18228_127 = 1'h1;
  assign T_18228_128 = T_16539;
  assign T_18228_129 = T_16562;
  assign T_18228_130 = 1'h1;
  assign T_18228_131 = 1'h1;
  assign T_18228_132 = 1'h1;
  assign T_18228_133 = 1'h1;
  assign T_18228_134 = 1'h1;
  assign T_18228_135 = 1'h1;
  assign T_18228_136 = 1'h1;
  assign T_18228_137 = 1'h1;
  assign T_18228_138 = 1'h1;
  assign T_18228_139 = 1'h1;
  assign T_18228_140 = 1'h1;
  assign T_18228_141 = 1'h1;
  assign T_18228_142 = 1'h1;
  assign T_18228_143 = 1'h1;
  assign T_18228_144 = 1'h1;
  assign T_18228_145 = 1'h1;
  assign T_18228_146 = 1'h1;
  assign T_18228_147 = 1'h1;
  assign T_18228_148 = 1'h1;
  assign T_18228_149 = 1'h1;
  assign T_18228_150 = 1'h1;
  assign T_18228_151 = 1'h1;
  assign T_18228_152 = 1'h1;
  assign T_18228_153 = 1'h1;
  assign T_18228_154 = 1'h1;
  assign T_18228_155 = 1'h1;
  assign T_18228_156 = 1'h1;
  assign T_18228_157 = 1'h1;
  assign T_18228_158 = 1'h1;
  assign T_18228_159 = 1'h1;
  assign T_18228_160 = 1'h1;
  assign T_18228_161 = 1'h1;
  assign T_18228_162 = 1'h1;
  assign T_18228_163 = 1'h1;
  assign T_18228_164 = 1'h1;
  assign T_18228_165 = 1'h1;
  assign T_18228_166 = 1'h1;
  assign T_18228_167 = 1'h1;
  assign T_18228_168 = 1'h1;
  assign T_18228_169 = 1'h1;
  assign T_18228_170 = 1'h1;
  assign T_18228_171 = 1'h1;
  assign T_18228_172 = 1'h1;
  assign T_18228_173 = 1'h1;
  assign T_18228_174 = 1'h1;
  assign T_18228_175 = 1'h1;
  assign T_18228_176 = 1'h1;
  assign T_18228_177 = 1'h1;
  assign T_18228_178 = 1'h1;
  assign T_18228_179 = 1'h1;
  assign T_18228_180 = 1'h1;
  assign T_18228_181 = 1'h1;
  assign T_18228_182 = 1'h1;
  assign T_18228_183 = 1'h1;
  assign T_18228_184 = 1'h1;
  assign T_18228_185 = 1'h1;
  assign T_18228_186 = 1'h1;
  assign T_18228_187 = 1'h1;
  assign T_18228_188 = 1'h1;
  assign T_18228_189 = 1'h1;
  assign T_18228_190 = 1'h1;
  assign T_18228_191 = 1'h1;
  assign T_18228_192 = 1'h1;
  assign T_18228_193 = 1'h1;
  assign T_18228_194 = 1'h1;
  assign T_18228_195 = 1'h1;
  assign T_18228_196 = 1'h1;
  assign T_18228_197 = 1'h1;
  assign T_18228_198 = 1'h1;
  assign T_18228_199 = 1'h1;
  assign T_18228_200 = 1'h1;
  assign T_18228_201 = 1'h1;
  assign T_18228_202 = 1'h1;
  assign T_18228_203 = 1'h1;
  assign T_18228_204 = 1'h1;
  assign T_18228_205 = 1'h1;
  assign T_18228_206 = 1'h1;
  assign T_18228_207 = 1'h1;
  assign T_18228_208 = 1'h1;
  assign T_18228_209 = 1'h1;
  assign T_18228_210 = 1'h1;
  assign T_18228_211 = 1'h1;
  assign T_18228_212 = 1'h1;
  assign T_18228_213 = 1'h1;
  assign T_18228_214 = 1'h1;
  assign T_18228_215 = 1'h1;
  assign T_18228_216 = 1'h1;
  assign T_18228_217 = 1'h1;
  assign T_18228_218 = 1'h1;
  assign T_18228_219 = 1'h1;
  assign T_18228_220 = 1'h1;
  assign T_18228_221 = 1'h1;
  assign T_18228_222 = 1'h1;
  assign T_18228_223 = 1'h1;
  assign T_18228_224 = 1'h1;
  assign T_18228_225 = 1'h1;
  assign T_18228_226 = 1'h1;
  assign T_18228_227 = 1'h1;
  assign T_18228_228 = 1'h1;
  assign T_18228_229 = 1'h1;
  assign T_18228_230 = 1'h1;
  assign T_18228_231 = 1'h1;
  assign T_18228_232 = 1'h1;
  assign T_18228_233 = 1'h1;
  assign T_18228_234 = 1'h1;
  assign T_18228_235 = 1'h1;
  assign T_18228_236 = 1'h1;
  assign T_18228_237 = 1'h1;
  assign T_18228_238 = 1'h1;
  assign T_18228_239 = 1'h1;
  assign T_18228_240 = 1'h1;
  assign T_18228_241 = 1'h1;
  assign T_18228_242 = 1'h1;
  assign T_18228_243 = 1'h1;
  assign T_18228_244 = 1'h1;
  assign T_18228_245 = 1'h1;
  assign T_18228_246 = 1'h1;
  assign T_18228_247 = 1'h1;
  assign T_18228_248 = 1'h1;
  assign T_18228_249 = 1'h1;
  assign T_18228_250 = 1'h1;
  assign T_18228_251 = 1'h1;
  assign T_18228_252 = 1'h1;
  assign T_18228_253 = 1'h1;
  assign T_18228_254 = 1'h1;
  assign T_18228_255 = 1'h1;
  assign T_18228_256 = T_4324_78;
  assign T_18228_257 = T_4324_63;
  assign T_18228_258 = 1'h1;
  assign T_18228_259 = 1'h1;
  assign T_18228_260 = 1'h1;
  assign T_18228_261 = 1'h1;
  assign T_18228_262 = 1'h1;
  assign T_18228_263 = 1'h1;
  assign T_18228_264 = 1'h1;
  assign T_18228_265 = 1'h1;
  assign T_18228_266 = 1'h1;
  assign T_18228_267 = 1'h1;
  assign T_18228_268 = 1'h1;
  assign T_18228_269 = 1'h1;
  assign T_18228_270 = 1'h1;
  assign T_18228_271 = 1'h1;
  assign T_18228_272 = 1'h1;
  assign T_18228_273 = 1'h1;
  assign T_18228_274 = 1'h1;
  assign T_18228_275 = 1'h1;
  assign T_18228_276 = 1'h1;
  assign T_18228_277 = 1'h1;
  assign T_18228_278 = 1'h1;
  assign T_18228_279 = 1'h1;
  assign T_18228_280 = 1'h1;
  assign T_18228_281 = 1'h1;
  assign T_18228_282 = 1'h1;
  assign T_18228_283 = 1'h1;
  assign T_18228_284 = 1'h1;
  assign T_18228_285 = 1'h1;
  assign T_18228_286 = 1'h1;
  assign T_18228_287 = 1'h1;
  assign T_18228_288 = 1'h1;
  assign T_18228_289 = 1'h1;
  assign T_18228_290 = 1'h1;
  assign T_18228_291 = 1'h1;
  assign T_18228_292 = 1'h1;
  assign T_18228_293 = 1'h1;
  assign T_18228_294 = 1'h1;
  assign T_18228_295 = 1'h1;
  assign T_18228_296 = 1'h1;
  assign T_18228_297 = 1'h1;
  assign T_18228_298 = 1'h1;
  assign T_18228_299 = 1'h1;
  assign T_18228_300 = 1'h1;
  assign T_18228_301 = 1'h1;
  assign T_18228_302 = 1'h1;
  assign T_18228_303 = 1'h1;
  assign T_18228_304 = 1'h1;
  assign T_18228_305 = 1'h1;
  assign T_18228_306 = 1'h1;
  assign T_18228_307 = 1'h1;
  assign T_18228_308 = 1'h1;
  assign T_18228_309 = 1'h1;
  assign T_18228_310 = 1'h1;
  assign T_18228_311 = 1'h1;
  assign T_18228_312 = 1'h1;
  assign T_18228_313 = 1'h1;
  assign T_18228_314 = 1'h1;
  assign T_18228_315 = 1'h1;
  assign T_18228_316 = 1'h1;
  assign T_18228_317 = 1'h1;
  assign T_18228_318 = 1'h1;
  assign T_18228_319 = 1'h1;
  assign T_18228_320 = 1'h1;
  assign T_18228_321 = 1'h1;
  assign T_18228_322 = 1'h1;
  assign T_18228_323 = 1'h1;
  assign T_18228_324 = 1'h1;
  assign T_18228_325 = 1'h1;
  assign T_18228_326 = 1'h1;
  assign T_18228_327 = 1'h1;
  assign T_18228_328 = 1'h1;
  assign T_18228_329 = 1'h1;
  assign T_18228_330 = 1'h1;
  assign T_18228_331 = 1'h1;
  assign T_18228_332 = 1'h1;
  assign T_18228_333 = 1'h1;
  assign T_18228_334 = 1'h1;
  assign T_18228_335 = 1'h1;
  assign T_18228_336 = 1'h1;
  assign T_18228_337 = 1'h1;
  assign T_18228_338 = 1'h1;
  assign T_18228_339 = 1'h1;
  assign T_18228_340 = 1'h1;
  assign T_18228_341 = 1'h1;
  assign T_18228_342 = 1'h1;
  assign T_18228_343 = 1'h1;
  assign T_18228_344 = 1'h1;
  assign T_18228_345 = 1'h1;
  assign T_18228_346 = 1'h1;
  assign T_18228_347 = 1'h1;
  assign T_18228_348 = 1'h1;
  assign T_18228_349 = 1'h1;
  assign T_18228_350 = 1'h1;
  assign T_18228_351 = 1'h1;
  assign T_18228_352 = 1'h1;
  assign T_18228_353 = 1'h1;
  assign T_18228_354 = 1'h1;
  assign T_18228_355 = 1'h1;
  assign T_18228_356 = 1'h1;
  assign T_18228_357 = 1'h1;
  assign T_18228_358 = 1'h1;
  assign T_18228_359 = 1'h1;
  assign T_18228_360 = 1'h1;
  assign T_18228_361 = 1'h1;
  assign T_18228_362 = 1'h1;
  assign T_18228_363 = 1'h1;
  assign T_18228_364 = 1'h1;
  assign T_18228_365 = 1'h1;
  assign T_18228_366 = 1'h1;
  assign T_18228_367 = 1'h1;
  assign T_18228_368 = 1'h1;
  assign T_18228_369 = 1'h1;
  assign T_18228_370 = 1'h1;
  assign T_18228_371 = 1'h1;
  assign T_18228_372 = 1'h1;
  assign T_18228_373 = 1'h1;
  assign T_18228_374 = 1'h1;
  assign T_18228_375 = 1'h1;
  assign T_18228_376 = 1'h1;
  assign T_18228_377 = 1'h1;
  assign T_18228_378 = 1'h1;
  assign T_18228_379 = 1'h1;
  assign T_18228_380 = 1'h1;
  assign T_18228_381 = 1'h1;
  assign T_18228_382 = 1'h1;
  assign T_18228_383 = 1'h1;
  assign T_18228_384 = 1'h1;
  assign T_18228_385 = 1'h1;
  assign T_18228_386 = 1'h1;
  assign T_18228_387 = 1'h1;
  assign T_18228_388 = 1'h1;
  assign T_18228_389 = 1'h1;
  assign T_18228_390 = 1'h1;
  assign T_18228_391 = 1'h1;
  assign T_18228_392 = 1'h1;
  assign T_18228_393 = 1'h1;
  assign T_18228_394 = 1'h1;
  assign T_18228_395 = 1'h1;
  assign T_18228_396 = 1'h1;
  assign T_18228_397 = 1'h1;
  assign T_18228_398 = 1'h1;
  assign T_18228_399 = 1'h1;
  assign T_18228_400 = 1'h1;
  assign T_18228_401 = 1'h1;
  assign T_18228_402 = 1'h1;
  assign T_18228_403 = 1'h1;
  assign T_18228_404 = 1'h1;
  assign T_18228_405 = 1'h1;
  assign T_18228_406 = 1'h1;
  assign T_18228_407 = 1'h1;
  assign T_18228_408 = 1'h1;
  assign T_18228_409 = 1'h1;
  assign T_18228_410 = 1'h1;
  assign T_18228_411 = 1'h1;
  assign T_18228_412 = 1'h1;
  assign T_18228_413 = 1'h1;
  assign T_18228_414 = 1'h1;
  assign T_18228_415 = 1'h1;
  assign T_18228_416 = 1'h1;
  assign T_18228_417 = 1'h1;
  assign T_18228_418 = 1'h1;
  assign T_18228_419 = 1'h1;
  assign T_18228_420 = 1'h1;
  assign T_18228_421 = 1'h1;
  assign T_18228_422 = 1'h1;
  assign T_18228_423 = 1'h1;
  assign T_18228_424 = 1'h1;
  assign T_18228_425 = 1'h1;
  assign T_18228_426 = 1'h1;
  assign T_18228_427 = 1'h1;
  assign T_18228_428 = 1'h1;
  assign T_18228_429 = 1'h1;
  assign T_18228_430 = 1'h1;
  assign T_18228_431 = 1'h1;
  assign T_18228_432 = 1'h1;
  assign T_18228_433 = 1'h1;
  assign T_18228_434 = 1'h1;
  assign T_18228_435 = 1'h1;
  assign T_18228_436 = 1'h1;
  assign T_18228_437 = 1'h1;
  assign T_18228_438 = 1'h1;
  assign T_18228_439 = 1'h1;
  assign T_18228_440 = 1'h1;
  assign T_18228_441 = 1'h1;
  assign T_18228_442 = 1'h1;
  assign T_18228_443 = 1'h1;
  assign T_18228_444 = 1'h1;
  assign T_18228_445 = 1'h1;
  assign T_18228_446 = 1'h1;
  assign T_18228_447 = 1'h1;
  assign T_18228_448 = 1'h1;
  assign T_18228_449 = 1'h1;
  assign T_18228_450 = 1'h1;
  assign T_18228_451 = 1'h1;
  assign T_18228_452 = 1'h1;
  assign T_18228_453 = 1'h1;
  assign T_18228_454 = 1'h1;
  assign T_18228_455 = 1'h1;
  assign T_18228_456 = 1'h1;
  assign T_18228_457 = 1'h1;
  assign T_18228_458 = 1'h1;
  assign T_18228_459 = 1'h1;
  assign T_18228_460 = 1'h1;
  assign T_18228_461 = 1'h1;
  assign T_18228_462 = 1'h1;
  assign T_18228_463 = 1'h1;
  assign T_18228_464 = 1'h1;
  assign T_18228_465 = 1'h1;
  assign T_18228_466 = 1'h1;
  assign T_18228_467 = 1'h1;
  assign T_18228_468 = 1'h1;
  assign T_18228_469 = 1'h1;
  assign T_18228_470 = 1'h1;
  assign T_18228_471 = 1'h1;
  assign T_18228_472 = 1'h1;
  assign T_18228_473 = 1'h1;
  assign T_18228_474 = 1'h1;
  assign T_18228_475 = 1'h1;
  assign T_18228_476 = 1'h1;
  assign T_18228_477 = 1'h1;
  assign T_18228_478 = 1'h1;
  assign T_18228_479 = 1'h1;
  assign T_18228_480 = 1'h1;
  assign T_18228_481 = 1'h1;
  assign T_18228_482 = 1'h1;
  assign T_18228_483 = 1'h1;
  assign T_18228_484 = 1'h1;
  assign T_18228_485 = 1'h1;
  assign T_18228_486 = 1'h1;
  assign T_18228_487 = 1'h1;
  assign T_18228_488 = 1'h1;
  assign T_18228_489 = 1'h1;
  assign T_18228_490 = 1'h1;
  assign T_18228_491 = 1'h1;
  assign T_18228_492 = 1'h1;
  assign T_18228_493 = 1'h1;
  assign T_18228_494 = 1'h1;
  assign T_18228_495 = 1'h1;
  assign T_18228_496 = 1'h1;
  assign T_18228_497 = 1'h1;
  assign T_18228_498 = 1'h1;
  assign T_18228_499 = 1'h1;
  assign T_18228_500 = 1'h1;
  assign T_18228_501 = 1'h1;
  assign T_18228_502 = 1'h1;
  assign T_18228_503 = 1'h1;
  assign T_18228_504 = 1'h1;
  assign T_18228_505 = 1'h1;
  assign T_18228_506 = 1'h1;
  assign T_18228_507 = 1'h1;
  assign T_18228_508 = 1'h1;
  assign T_18228_509 = 1'h1;
  assign T_18228_510 = 1'h1;
  assign T_18228_511 = 1'h1;
  assign T_18989 = T_4329_31 & T_4329_30;
  assign T_18990 = T_18989 & T_4329_29;
  assign T_18991 = T_18990 & T_4329_28;
  assign T_18992 = T_18991 & T_4329_27;
  assign T_18993 = T_18992 & T_4329_26;
  assign T_18994 = T_18993 & T_4329_25;
  assign T_18995 = T_18994 & T_4329_24;
  assign T_18996 = T_18995 & T_4329_23;
  assign T_18997 = T_18996 & T_4329_22;
  assign T_18998 = T_18997 & T_4329_21;
  assign T_18999 = T_18998 & T_4329_20;
  assign T_19000 = T_18999 & T_4329_19;
  assign T_19001 = T_19000 & T_4329_18;
  assign T_19002 = T_19001 & T_4329_17;
  assign T_19003 = T_19002 & T_4329_16;
  assign T_19004 = T_19003 & T_4329_15;
  assign T_19005 = T_19004 & T_4329_14;
  assign T_19006 = T_19005 & T_4329_13;
  assign T_19007 = T_19006 & T_4329_12;
  assign T_19008 = T_19007 & T_4329_11;
  assign T_19009 = T_19008 & T_4329_10;
  assign T_19010 = T_19009 & T_4329_9;
  assign T_19011 = T_19010 & T_4329_8;
  assign T_19012 = T_19011 & T_4329_7;
  assign T_19013 = T_19012 & T_4329_6;
  assign T_19014 = T_19013 & T_4329_5;
  assign T_19015 = T_19014 & T_4329_4;
  assign T_19016 = T_19015 & T_4329_3;
  assign T_19017 = T_19016 & T_4329_2;
  assign T_19018 = T_19017 & T_4329_1;
  assign T_19019 = T_19018 & T_4329_0;
  assign T_19024 = T_4329_140 & T_4329_139;
  assign T_19025 = T_19024 & T_4329_138;
  assign T_19026 = T_19025 & T_4329_137;
  assign T_19027 = T_19026 & T_4329_136;
  assign T_19028 = T_19027 & T_4329_135;
  assign T_19029 = T_19028 & T_4329_134;
  assign T_19030 = T_19029 & T_4329_133;
  assign T_19031 = T_19030 & T_4329_132;
  assign T_19032 = T_19031 & T_4329_131;
  assign T_19033 = T_19032 & T_4329_130;
  assign T_19034 = T_19033 & T_4329_129;
  assign T_19035 = T_19034 & T_4329_128;
  assign T_19036 = T_19035 & T_4329_127;
  assign T_19037 = T_19036 & T_4329_126;
  assign T_19038 = T_19037 & T_4329_125;
  assign T_19039 = T_19038 & T_4329_124;
  assign T_19040 = T_19039 & T_4329_123;
  assign T_19041 = T_19040 & T_4329_122;
  assign T_19042 = T_19041 & T_4329_121;
  assign T_19233 = T_4329_110 & T_4329_109;
  assign T_19234 = T_19233 & T_4329_108;
  assign T_19235 = T_19234 & T_4329_107;
  assign T_19236 = T_19235 & T_4329_106;
  assign T_19237 = T_19236 & T_4329_105;
  assign T_19238 = T_19237 & T_4329_104;
  assign T_19239 = T_19238 & T_4329_103;
  assign T_19240 = T_19239 & T_4329_102;
  assign T_19241 = T_19240 & T_4329_101;
  assign T_19242 = T_19241 & T_4329_100;
  assign T_19243 = T_19242 & T_4329_99;
  assign T_19244 = T_19243 & T_4329_98;
  assign T_19245 = T_19244 & T_4329_97;
  assign T_19246 = T_19245 & T_4329_96;
  assign T_19247 = T_19246 & T_4329_95;
  assign T_19248 = T_19247 & T_4329_94;
  assign T_19249 = T_19248 & T_4329_93;
  assign T_19250 = T_19249 & T_4329_92;
  assign T_19251 = T_19250 & T_4329_91;
  assign T_19252 = T_19251 & T_4329_90;
  assign T_19253 = T_19252 & T_4329_89;
  assign T_19254 = T_19253 & T_4329_88;
  assign T_19255 = T_19254 & T_4329_87;
  assign T_19256 = T_19255 & T_4329_86;
  assign T_19257 = T_19256 & T_4329_85;
  assign T_19258 = T_19257 & T_4329_84;
  assign T_19259 = T_19258 & T_4329_83;
  assign T_19260 = T_19259 & T_4329_82;
  assign T_19261 = T_19260 & T_4329_81;
  assign T_19262 = T_19261 & T_4329_80;
  assign T_19263 = T_19262 & T_4329_79;
  assign T_19268 = T_4329_60 & T_4329_59;
  assign T_19269 = T_19268 & T_4329_58;
  assign T_19270 = T_19269 & T_4329_57;
  assign T_19271 = T_19270 & T_4329_56;
  assign T_19272 = T_19271 & T_4329_55;
  assign T_19273 = T_19272 & T_4329_54;
  assign T_19274 = T_19273 & T_4329_53;
  assign T_19275 = T_19274 & T_4329_52;
  assign T_19276 = T_19275 & T_4329_51;
  assign T_19277 = T_19276 & T_4329_50;
  assign T_19278 = T_19277 & T_4329_49;
  assign T_19279 = T_19278 & T_4329_48;
  assign T_19280 = T_19279 & T_4329_47;
  assign T_19281 = T_19280 & T_4329_46;
  assign T_19282 = T_19281 & T_4329_45;
  assign T_19283 = T_19282 & T_4329_44;
  assign T_19284 = T_19283 & T_4329_43;
  assign T_19285 = T_19284 & T_4329_42;
  assign T_19286 = T_19285 & T_4329_41;
  assign T_20952_0 = T_4329_32;
  assign T_20952_1 = T_4329_64;
  assign T_20952_2 = T_4329_73;
  assign T_20952_3 = T_4329_118;
  assign T_20952_4 = T_4329_155;
  assign T_20952_5 = T_4329_33;
  assign T_20952_6 = T_4329_65;
  assign T_20952_7 = T_4329_116;
  assign T_20952_8 = T_4329_150;
  assign T_20952_9 = T_4329_70;
  assign T_20952_10 = T_4329_34;
  assign T_20952_11 = T_4329_145;
  assign T_20952_12 = T_4329_114;
  assign T_20952_13 = T_4329_71;
  assign T_20952_14 = T_4329_39;
  assign T_20952_15 = T_4329_157;
  assign T_20952_16 = T_4329_143;
  assign T_20952_17 = T_4329_77;
  assign T_20952_18 = T_4329_141;
  assign T_20952_19 = T_4329_154;
  assign T_20952_20 = T_4329_40;
  assign T_20952_21 = T_4329_68;
  assign T_20952_22 = T_4329_111;
  assign T_20952_23 = T_4329_149;
  assign T_20952_24 = T_4329_36;
  assign T_20952_25 = T_4329_38;
  assign T_20952_26 = T_4329_148;
  assign T_20952_27 = T_4329_113;
  assign T_20952_28 = T_4329_66;
  assign T_20952_29 = T_4329_62;
  assign T_20952_30 = T_4329_152;
  assign T_20952_31 = T_4329_144;
  assign T_20952_32 = T_4329_74;
  assign T_20952_33 = T_4329_69;
  assign T_20952_34 = T_4329_75;
  assign T_20952_35 = T_4329_119;
  assign T_20952_36 = T_4329_151;
  assign T_20952_37 = T_4329_37;
  assign T_20952_38 = T_4329_67;
  assign T_20952_39 = T_4329_117;
  assign T_20952_40 = T_4329_147;
  assign T_20952_41 = T_4329_72;
  assign T_20952_42 = T_4329_35;
  assign T_20952_43 = T_4329_146;
  assign T_20952_44 = T_4329_112;
  assign T_20952_45 = T_4329_76;
  assign T_20952_46 = T_4329_61;
  assign T_20952_47 = T_4329_156;
  assign T_20952_48 = T_4329_120;
  assign T_20952_49 = T_4329_115;
  assign T_20952_50 = T_4329_142;
  assign T_20952_51 = T_4329_153;
  assign T_20952_52 = 1'h1;
  assign T_20952_53 = 1'h1;
  assign T_20952_54 = 1'h1;
  assign T_20952_55 = 1'h1;
  assign T_20952_56 = 1'h1;
  assign T_20952_57 = 1'h1;
  assign T_20952_58 = 1'h1;
  assign T_20952_59 = 1'h1;
  assign T_20952_60 = 1'h1;
  assign T_20952_61 = 1'h1;
  assign T_20952_62 = 1'h1;
  assign T_20952_63 = 1'h1;
  assign T_20952_64 = T_19019;
  assign T_20952_65 = T_19042;
  assign T_20952_66 = 1'h1;
  assign T_20952_67 = 1'h1;
  assign T_20952_68 = 1'h1;
  assign T_20952_69 = 1'h1;
  assign T_20952_70 = 1'h1;
  assign T_20952_71 = 1'h1;
  assign T_20952_72 = 1'h1;
  assign T_20952_73 = 1'h1;
  assign T_20952_74 = 1'h1;
  assign T_20952_75 = 1'h1;
  assign T_20952_76 = 1'h1;
  assign T_20952_77 = 1'h1;
  assign T_20952_78 = 1'h1;
  assign T_20952_79 = 1'h1;
  assign T_20952_80 = 1'h1;
  assign T_20952_81 = 1'h1;
  assign T_20952_82 = 1'h1;
  assign T_20952_83 = 1'h1;
  assign T_20952_84 = 1'h1;
  assign T_20952_85 = 1'h1;
  assign T_20952_86 = 1'h1;
  assign T_20952_87 = 1'h1;
  assign T_20952_88 = 1'h1;
  assign T_20952_89 = 1'h1;
  assign T_20952_90 = 1'h1;
  assign T_20952_91 = 1'h1;
  assign T_20952_92 = 1'h1;
  assign T_20952_93 = 1'h1;
  assign T_20952_94 = 1'h1;
  assign T_20952_95 = 1'h1;
  assign T_20952_96 = 1'h1;
  assign T_20952_97 = 1'h1;
  assign T_20952_98 = 1'h1;
  assign T_20952_99 = 1'h1;
  assign T_20952_100 = 1'h1;
  assign T_20952_101 = 1'h1;
  assign T_20952_102 = 1'h1;
  assign T_20952_103 = 1'h1;
  assign T_20952_104 = 1'h1;
  assign T_20952_105 = 1'h1;
  assign T_20952_106 = 1'h1;
  assign T_20952_107 = 1'h1;
  assign T_20952_108 = 1'h1;
  assign T_20952_109 = 1'h1;
  assign T_20952_110 = 1'h1;
  assign T_20952_111 = 1'h1;
  assign T_20952_112 = 1'h1;
  assign T_20952_113 = 1'h1;
  assign T_20952_114 = 1'h1;
  assign T_20952_115 = 1'h1;
  assign T_20952_116 = 1'h1;
  assign T_20952_117 = 1'h1;
  assign T_20952_118 = 1'h1;
  assign T_20952_119 = 1'h1;
  assign T_20952_120 = 1'h1;
  assign T_20952_121 = 1'h1;
  assign T_20952_122 = 1'h1;
  assign T_20952_123 = 1'h1;
  assign T_20952_124 = 1'h1;
  assign T_20952_125 = 1'h1;
  assign T_20952_126 = 1'h1;
  assign T_20952_127 = 1'h1;
  assign T_20952_128 = T_19263;
  assign T_20952_129 = T_19286;
  assign T_20952_130 = 1'h1;
  assign T_20952_131 = 1'h1;
  assign T_20952_132 = 1'h1;
  assign T_20952_133 = 1'h1;
  assign T_20952_134 = 1'h1;
  assign T_20952_135 = 1'h1;
  assign T_20952_136 = 1'h1;
  assign T_20952_137 = 1'h1;
  assign T_20952_138 = 1'h1;
  assign T_20952_139 = 1'h1;
  assign T_20952_140 = 1'h1;
  assign T_20952_141 = 1'h1;
  assign T_20952_142 = 1'h1;
  assign T_20952_143 = 1'h1;
  assign T_20952_144 = 1'h1;
  assign T_20952_145 = 1'h1;
  assign T_20952_146 = 1'h1;
  assign T_20952_147 = 1'h1;
  assign T_20952_148 = 1'h1;
  assign T_20952_149 = 1'h1;
  assign T_20952_150 = 1'h1;
  assign T_20952_151 = 1'h1;
  assign T_20952_152 = 1'h1;
  assign T_20952_153 = 1'h1;
  assign T_20952_154 = 1'h1;
  assign T_20952_155 = 1'h1;
  assign T_20952_156 = 1'h1;
  assign T_20952_157 = 1'h1;
  assign T_20952_158 = 1'h1;
  assign T_20952_159 = 1'h1;
  assign T_20952_160 = 1'h1;
  assign T_20952_161 = 1'h1;
  assign T_20952_162 = 1'h1;
  assign T_20952_163 = 1'h1;
  assign T_20952_164 = 1'h1;
  assign T_20952_165 = 1'h1;
  assign T_20952_166 = 1'h1;
  assign T_20952_167 = 1'h1;
  assign T_20952_168 = 1'h1;
  assign T_20952_169 = 1'h1;
  assign T_20952_170 = 1'h1;
  assign T_20952_171 = 1'h1;
  assign T_20952_172 = 1'h1;
  assign T_20952_173 = 1'h1;
  assign T_20952_174 = 1'h1;
  assign T_20952_175 = 1'h1;
  assign T_20952_176 = 1'h1;
  assign T_20952_177 = 1'h1;
  assign T_20952_178 = 1'h1;
  assign T_20952_179 = 1'h1;
  assign T_20952_180 = 1'h1;
  assign T_20952_181 = 1'h1;
  assign T_20952_182 = 1'h1;
  assign T_20952_183 = 1'h1;
  assign T_20952_184 = 1'h1;
  assign T_20952_185 = 1'h1;
  assign T_20952_186 = 1'h1;
  assign T_20952_187 = 1'h1;
  assign T_20952_188 = 1'h1;
  assign T_20952_189 = 1'h1;
  assign T_20952_190 = 1'h1;
  assign T_20952_191 = 1'h1;
  assign T_20952_192 = 1'h1;
  assign T_20952_193 = 1'h1;
  assign T_20952_194 = 1'h1;
  assign T_20952_195 = 1'h1;
  assign T_20952_196 = 1'h1;
  assign T_20952_197 = 1'h1;
  assign T_20952_198 = 1'h1;
  assign T_20952_199 = 1'h1;
  assign T_20952_200 = 1'h1;
  assign T_20952_201 = 1'h1;
  assign T_20952_202 = 1'h1;
  assign T_20952_203 = 1'h1;
  assign T_20952_204 = 1'h1;
  assign T_20952_205 = 1'h1;
  assign T_20952_206 = 1'h1;
  assign T_20952_207 = 1'h1;
  assign T_20952_208 = 1'h1;
  assign T_20952_209 = 1'h1;
  assign T_20952_210 = 1'h1;
  assign T_20952_211 = 1'h1;
  assign T_20952_212 = 1'h1;
  assign T_20952_213 = 1'h1;
  assign T_20952_214 = 1'h1;
  assign T_20952_215 = 1'h1;
  assign T_20952_216 = 1'h1;
  assign T_20952_217 = 1'h1;
  assign T_20952_218 = 1'h1;
  assign T_20952_219 = 1'h1;
  assign T_20952_220 = 1'h1;
  assign T_20952_221 = 1'h1;
  assign T_20952_222 = 1'h1;
  assign T_20952_223 = 1'h1;
  assign T_20952_224 = 1'h1;
  assign T_20952_225 = 1'h1;
  assign T_20952_226 = 1'h1;
  assign T_20952_227 = 1'h1;
  assign T_20952_228 = 1'h1;
  assign T_20952_229 = 1'h1;
  assign T_20952_230 = 1'h1;
  assign T_20952_231 = 1'h1;
  assign T_20952_232 = 1'h1;
  assign T_20952_233 = 1'h1;
  assign T_20952_234 = 1'h1;
  assign T_20952_235 = 1'h1;
  assign T_20952_236 = 1'h1;
  assign T_20952_237 = 1'h1;
  assign T_20952_238 = 1'h1;
  assign T_20952_239 = 1'h1;
  assign T_20952_240 = 1'h1;
  assign T_20952_241 = 1'h1;
  assign T_20952_242 = 1'h1;
  assign T_20952_243 = 1'h1;
  assign T_20952_244 = 1'h1;
  assign T_20952_245 = 1'h1;
  assign T_20952_246 = 1'h1;
  assign T_20952_247 = 1'h1;
  assign T_20952_248 = 1'h1;
  assign T_20952_249 = 1'h1;
  assign T_20952_250 = 1'h1;
  assign T_20952_251 = 1'h1;
  assign T_20952_252 = 1'h1;
  assign T_20952_253 = 1'h1;
  assign T_20952_254 = 1'h1;
  assign T_20952_255 = 1'h1;
  assign T_20952_256 = T_4329_78;
  assign T_20952_257 = T_4329_63;
  assign T_20952_258 = 1'h1;
  assign T_20952_259 = 1'h1;
  assign T_20952_260 = 1'h1;
  assign T_20952_261 = 1'h1;
  assign T_20952_262 = 1'h1;
  assign T_20952_263 = 1'h1;
  assign T_20952_264 = 1'h1;
  assign T_20952_265 = 1'h1;
  assign T_20952_266 = 1'h1;
  assign T_20952_267 = 1'h1;
  assign T_20952_268 = 1'h1;
  assign T_20952_269 = 1'h1;
  assign T_20952_270 = 1'h1;
  assign T_20952_271 = 1'h1;
  assign T_20952_272 = 1'h1;
  assign T_20952_273 = 1'h1;
  assign T_20952_274 = 1'h1;
  assign T_20952_275 = 1'h1;
  assign T_20952_276 = 1'h1;
  assign T_20952_277 = 1'h1;
  assign T_20952_278 = 1'h1;
  assign T_20952_279 = 1'h1;
  assign T_20952_280 = 1'h1;
  assign T_20952_281 = 1'h1;
  assign T_20952_282 = 1'h1;
  assign T_20952_283 = 1'h1;
  assign T_20952_284 = 1'h1;
  assign T_20952_285 = 1'h1;
  assign T_20952_286 = 1'h1;
  assign T_20952_287 = 1'h1;
  assign T_20952_288 = 1'h1;
  assign T_20952_289 = 1'h1;
  assign T_20952_290 = 1'h1;
  assign T_20952_291 = 1'h1;
  assign T_20952_292 = 1'h1;
  assign T_20952_293 = 1'h1;
  assign T_20952_294 = 1'h1;
  assign T_20952_295 = 1'h1;
  assign T_20952_296 = 1'h1;
  assign T_20952_297 = 1'h1;
  assign T_20952_298 = 1'h1;
  assign T_20952_299 = 1'h1;
  assign T_20952_300 = 1'h1;
  assign T_20952_301 = 1'h1;
  assign T_20952_302 = 1'h1;
  assign T_20952_303 = 1'h1;
  assign T_20952_304 = 1'h1;
  assign T_20952_305 = 1'h1;
  assign T_20952_306 = 1'h1;
  assign T_20952_307 = 1'h1;
  assign T_20952_308 = 1'h1;
  assign T_20952_309 = 1'h1;
  assign T_20952_310 = 1'h1;
  assign T_20952_311 = 1'h1;
  assign T_20952_312 = 1'h1;
  assign T_20952_313 = 1'h1;
  assign T_20952_314 = 1'h1;
  assign T_20952_315 = 1'h1;
  assign T_20952_316 = 1'h1;
  assign T_20952_317 = 1'h1;
  assign T_20952_318 = 1'h1;
  assign T_20952_319 = 1'h1;
  assign T_20952_320 = 1'h1;
  assign T_20952_321 = 1'h1;
  assign T_20952_322 = 1'h1;
  assign T_20952_323 = 1'h1;
  assign T_20952_324 = 1'h1;
  assign T_20952_325 = 1'h1;
  assign T_20952_326 = 1'h1;
  assign T_20952_327 = 1'h1;
  assign T_20952_328 = 1'h1;
  assign T_20952_329 = 1'h1;
  assign T_20952_330 = 1'h1;
  assign T_20952_331 = 1'h1;
  assign T_20952_332 = 1'h1;
  assign T_20952_333 = 1'h1;
  assign T_20952_334 = 1'h1;
  assign T_20952_335 = 1'h1;
  assign T_20952_336 = 1'h1;
  assign T_20952_337 = 1'h1;
  assign T_20952_338 = 1'h1;
  assign T_20952_339 = 1'h1;
  assign T_20952_340 = 1'h1;
  assign T_20952_341 = 1'h1;
  assign T_20952_342 = 1'h1;
  assign T_20952_343 = 1'h1;
  assign T_20952_344 = 1'h1;
  assign T_20952_345 = 1'h1;
  assign T_20952_346 = 1'h1;
  assign T_20952_347 = 1'h1;
  assign T_20952_348 = 1'h1;
  assign T_20952_349 = 1'h1;
  assign T_20952_350 = 1'h1;
  assign T_20952_351 = 1'h1;
  assign T_20952_352 = 1'h1;
  assign T_20952_353 = 1'h1;
  assign T_20952_354 = 1'h1;
  assign T_20952_355 = 1'h1;
  assign T_20952_356 = 1'h1;
  assign T_20952_357 = 1'h1;
  assign T_20952_358 = 1'h1;
  assign T_20952_359 = 1'h1;
  assign T_20952_360 = 1'h1;
  assign T_20952_361 = 1'h1;
  assign T_20952_362 = 1'h1;
  assign T_20952_363 = 1'h1;
  assign T_20952_364 = 1'h1;
  assign T_20952_365 = 1'h1;
  assign T_20952_366 = 1'h1;
  assign T_20952_367 = 1'h1;
  assign T_20952_368 = 1'h1;
  assign T_20952_369 = 1'h1;
  assign T_20952_370 = 1'h1;
  assign T_20952_371 = 1'h1;
  assign T_20952_372 = 1'h1;
  assign T_20952_373 = 1'h1;
  assign T_20952_374 = 1'h1;
  assign T_20952_375 = 1'h1;
  assign T_20952_376 = 1'h1;
  assign T_20952_377 = 1'h1;
  assign T_20952_378 = 1'h1;
  assign T_20952_379 = 1'h1;
  assign T_20952_380 = 1'h1;
  assign T_20952_381 = 1'h1;
  assign T_20952_382 = 1'h1;
  assign T_20952_383 = 1'h1;
  assign T_20952_384 = 1'h1;
  assign T_20952_385 = 1'h1;
  assign T_20952_386 = 1'h1;
  assign T_20952_387 = 1'h1;
  assign T_20952_388 = 1'h1;
  assign T_20952_389 = 1'h1;
  assign T_20952_390 = 1'h1;
  assign T_20952_391 = 1'h1;
  assign T_20952_392 = 1'h1;
  assign T_20952_393 = 1'h1;
  assign T_20952_394 = 1'h1;
  assign T_20952_395 = 1'h1;
  assign T_20952_396 = 1'h1;
  assign T_20952_397 = 1'h1;
  assign T_20952_398 = 1'h1;
  assign T_20952_399 = 1'h1;
  assign T_20952_400 = 1'h1;
  assign T_20952_401 = 1'h1;
  assign T_20952_402 = 1'h1;
  assign T_20952_403 = 1'h1;
  assign T_20952_404 = 1'h1;
  assign T_20952_405 = 1'h1;
  assign T_20952_406 = 1'h1;
  assign T_20952_407 = 1'h1;
  assign T_20952_408 = 1'h1;
  assign T_20952_409 = 1'h1;
  assign T_20952_410 = 1'h1;
  assign T_20952_411 = 1'h1;
  assign T_20952_412 = 1'h1;
  assign T_20952_413 = 1'h1;
  assign T_20952_414 = 1'h1;
  assign T_20952_415 = 1'h1;
  assign T_20952_416 = 1'h1;
  assign T_20952_417 = 1'h1;
  assign T_20952_418 = 1'h1;
  assign T_20952_419 = 1'h1;
  assign T_20952_420 = 1'h1;
  assign T_20952_421 = 1'h1;
  assign T_20952_422 = 1'h1;
  assign T_20952_423 = 1'h1;
  assign T_20952_424 = 1'h1;
  assign T_20952_425 = 1'h1;
  assign T_20952_426 = 1'h1;
  assign T_20952_427 = 1'h1;
  assign T_20952_428 = 1'h1;
  assign T_20952_429 = 1'h1;
  assign T_20952_430 = 1'h1;
  assign T_20952_431 = 1'h1;
  assign T_20952_432 = 1'h1;
  assign T_20952_433 = 1'h1;
  assign T_20952_434 = 1'h1;
  assign T_20952_435 = 1'h1;
  assign T_20952_436 = 1'h1;
  assign T_20952_437 = 1'h1;
  assign T_20952_438 = 1'h1;
  assign T_20952_439 = 1'h1;
  assign T_20952_440 = 1'h1;
  assign T_20952_441 = 1'h1;
  assign T_20952_442 = 1'h1;
  assign T_20952_443 = 1'h1;
  assign T_20952_444 = 1'h1;
  assign T_20952_445 = 1'h1;
  assign T_20952_446 = 1'h1;
  assign T_20952_447 = 1'h1;
  assign T_20952_448 = 1'h1;
  assign T_20952_449 = 1'h1;
  assign T_20952_450 = 1'h1;
  assign T_20952_451 = 1'h1;
  assign T_20952_452 = 1'h1;
  assign T_20952_453 = 1'h1;
  assign T_20952_454 = 1'h1;
  assign T_20952_455 = 1'h1;
  assign T_20952_456 = 1'h1;
  assign T_20952_457 = 1'h1;
  assign T_20952_458 = 1'h1;
  assign T_20952_459 = 1'h1;
  assign T_20952_460 = 1'h1;
  assign T_20952_461 = 1'h1;
  assign T_20952_462 = 1'h1;
  assign T_20952_463 = 1'h1;
  assign T_20952_464 = 1'h1;
  assign T_20952_465 = 1'h1;
  assign T_20952_466 = 1'h1;
  assign T_20952_467 = 1'h1;
  assign T_20952_468 = 1'h1;
  assign T_20952_469 = 1'h1;
  assign T_20952_470 = 1'h1;
  assign T_20952_471 = 1'h1;
  assign T_20952_472 = 1'h1;
  assign T_20952_473 = 1'h1;
  assign T_20952_474 = 1'h1;
  assign T_20952_475 = 1'h1;
  assign T_20952_476 = 1'h1;
  assign T_20952_477 = 1'h1;
  assign T_20952_478 = 1'h1;
  assign T_20952_479 = 1'h1;
  assign T_20952_480 = 1'h1;
  assign T_20952_481 = 1'h1;
  assign T_20952_482 = 1'h1;
  assign T_20952_483 = 1'h1;
  assign T_20952_484 = 1'h1;
  assign T_20952_485 = 1'h1;
  assign T_20952_486 = 1'h1;
  assign T_20952_487 = 1'h1;
  assign T_20952_488 = 1'h1;
  assign T_20952_489 = 1'h1;
  assign T_20952_490 = 1'h1;
  assign T_20952_491 = 1'h1;
  assign T_20952_492 = 1'h1;
  assign T_20952_493 = 1'h1;
  assign T_20952_494 = 1'h1;
  assign T_20952_495 = 1'h1;
  assign T_20952_496 = 1'h1;
  assign T_20952_497 = 1'h1;
  assign T_20952_498 = 1'h1;
  assign T_20952_499 = 1'h1;
  assign T_20952_500 = 1'h1;
  assign T_20952_501 = 1'h1;
  assign T_20952_502 = 1'h1;
  assign T_20952_503 = 1'h1;
  assign T_20952_504 = 1'h1;
  assign T_20952_505 = 1'h1;
  assign T_20952_506 = 1'h1;
  assign T_20952_507 = 1'h1;
  assign T_20952_508 = 1'h1;
  assign T_20952_509 = 1'h1;
  assign T_20952_510 = 1'h1;
  assign T_20952_511 = 1'h1;
  assign T_21713 = T_4334_31 & T_4334_30;
  assign T_21714 = T_21713 & T_4334_29;
  assign T_21715 = T_21714 & T_4334_28;
  assign T_21716 = T_21715 & T_4334_27;
  assign T_21717 = T_21716 & T_4334_26;
  assign T_21718 = T_21717 & T_4334_25;
  assign T_21719 = T_21718 & T_4334_24;
  assign T_21720 = T_21719 & T_4334_23;
  assign T_21721 = T_21720 & T_4334_22;
  assign T_21722 = T_21721 & T_4334_21;
  assign T_21723 = T_21722 & T_4334_20;
  assign T_21724 = T_21723 & T_4334_19;
  assign T_21725 = T_21724 & T_4334_18;
  assign T_21726 = T_21725 & T_4334_17;
  assign T_21727 = T_21726 & T_4334_16;
  assign T_21728 = T_21727 & T_4334_15;
  assign T_21729 = T_21728 & T_4334_14;
  assign T_21730 = T_21729 & T_4334_13;
  assign T_21731 = T_21730 & T_4334_12;
  assign T_21732 = T_21731 & T_4334_11;
  assign T_21733 = T_21732 & T_4334_10;
  assign T_21734 = T_21733 & T_4334_9;
  assign T_21735 = T_21734 & T_4334_8;
  assign T_21736 = T_21735 & T_4334_7;
  assign T_21737 = T_21736 & T_4334_6;
  assign T_21738 = T_21737 & T_4334_5;
  assign T_21739 = T_21738 & T_4334_4;
  assign T_21740 = T_21739 & T_4334_3;
  assign T_21741 = T_21740 & T_4334_2;
  assign T_21742 = T_21741 & T_4334_1;
  assign T_21743 = T_21742 & T_4334_0;
  assign T_21748 = T_4334_140 & T_4334_139;
  assign T_21749 = T_21748 & T_4334_138;
  assign T_21750 = T_21749 & T_4334_137;
  assign T_21751 = T_21750 & T_4334_136;
  assign T_21752 = T_21751 & T_4334_135;
  assign T_21753 = T_21752 & T_4334_134;
  assign T_21754 = T_21753 & T_4334_133;
  assign T_21755 = T_21754 & T_4334_132;
  assign T_21756 = T_21755 & T_4334_131;
  assign T_21757 = T_21756 & T_4334_130;
  assign T_21758 = T_21757 & T_4334_129;
  assign T_21759 = T_21758 & T_4334_128;
  assign T_21760 = T_21759 & T_4334_127;
  assign T_21761 = T_21760 & T_4334_126;
  assign T_21762 = T_21761 & T_4334_125;
  assign T_21763 = T_21762 & T_4334_124;
  assign T_21764 = T_21763 & T_4334_123;
  assign T_21765 = T_21764 & T_4334_122;
  assign T_21766 = T_21765 & T_4334_121;
  assign T_21957 = T_4334_110 & T_4334_109;
  assign T_21958 = T_21957 & T_4334_108;
  assign T_21959 = T_21958 & T_4334_107;
  assign T_21960 = T_21959 & T_4334_106;
  assign T_21961 = T_21960 & T_4334_105;
  assign T_21962 = T_21961 & T_4334_104;
  assign T_21963 = T_21962 & T_4334_103;
  assign T_21964 = T_21963 & T_4334_102;
  assign T_21965 = T_21964 & T_4334_101;
  assign T_21966 = T_21965 & T_4334_100;
  assign T_21967 = T_21966 & T_4334_99;
  assign T_21968 = T_21967 & T_4334_98;
  assign T_21969 = T_21968 & T_4334_97;
  assign T_21970 = T_21969 & T_4334_96;
  assign T_21971 = T_21970 & T_4334_95;
  assign T_21972 = T_21971 & T_4334_94;
  assign T_21973 = T_21972 & T_4334_93;
  assign T_21974 = T_21973 & T_4334_92;
  assign T_21975 = T_21974 & T_4334_91;
  assign T_21976 = T_21975 & T_4334_90;
  assign T_21977 = T_21976 & T_4334_89;
  assign T_21978 = T_21977 & T_4334_88;
  assign T_21979 = T_21978 & T_4334_87;
  assign T_21980 = T_21979 & T_4334_86;
  assign T_21981 = T_21980 & T_4334_85;
  assign T_21982 = T_21981 & T_4334_84;
  assign T_21983 = T_21982 & T_4334_83;
  assign T_21984 = T_21983 & T_4334_82;
  assign T_21985 = T_21984 & T_4334_81;
  assign T_21986 = T_21985 & T_4334_80;
  assign T_21987 = T_21986 & T_4334_79;
  assign T_21992 = T_4334_60 & T_4334_59;
  assign T_21993 = T_21992 & T_4334_58;
  assign T_21994 = T_21993 & T_4334_57;
  assign T_21995 = T_21994 & T_4334_56;
  assign T_21996 = T_21995 & T_4334_55;
  assign T_21997 = T_21996 & T_4334_54;
  assign T_21998 = T_21997 & T_4334_53;
  assign T_21999 = T_21998 & T_4334_52;
  assign T_22000 = T_21999 & T_4334_51;
  assign T_22001 = T_22000 & T_4334_50;
  assign T_22002 = T_22001 & T_4334_49;
  assign T_22003 = T_22002 & T_4334_48;
  assign T_22004 = T_22003 & T_4334_47;
  assign T_22005 = T_22004 & T_4334_46;
  assign T_22006 = T_22005 & T_4334_45;
  assign T_22007 = T_22006 & T_4334_44;
  assign T_22008 = T_22007 & T_4334_43;
  assign T_22009 = T_22008 & T_4334_42;
  assign T_22010 = T_22009 & T_4334_41;
  assign T_23676_0 = T_4334_32;
  assign T_23676_1 = T_4334_64;
  assign T_23676_2 = T_4334_73;
  assign T_23676_3 = T_4334_118;
  assign T_23676_4 = T_4334_155;
  assign T_23676_5 = T_4334_33;
  assign T_23676_6 = T_4334_65;
  assign T_23676_7 = T_4334_116;
  assign T_23676_8 = T_4334_150;
  assign T_23676_9 = T_4334_70;
  assign T_23676_10 = T_4334_34;
  assign T_23676_11 = T_4334_145;
  assign T_23676_12 = T_4334_114;
  assign T_23676_13 = T_4334_71;
  assign T_23676_14 = T_4334_39;
  assign T_23676_15 = T_4334_157;
  assign T_23676_16 = T_4334_143;
  assign T_23676_17 = T_4334_77;
  assign T_23676_18 = T_4334_141;
  assign T_23676_19 = T_4334_154;
  assign T_23676_20 = T_4334_40;
  assign T_23676_21 = T_4334_68;
  assign T_23676_22 = T_4334_111;
  assign T_23676_23 = T_4334_149;
  assign T_23676_24 = T_4334_36;
  assign T_23676_25 = T_4334_38;
  assign T_23676_26 = T_4334_148;
  assign T_23676_27 = T_4334_113;
  assign T_23676_28 = T_4334_66;
  assign T_23676_29 = T_4334_62;
  assign T_23676_30 = T_4334_152;
  assign T_23676_31 = T_4334_144;
  assign T_23676_32 = T_4334_74;
  assign T_23676_33 = T_4334_69;
  assign T_23676_34 = T_4334_75;
  assign T_23676_35 = T_4334_119;
  assign T_23676_36 = T_4334_151;
  assign T_23676_37 = T_4334_37;
  assign T_23676_38 = T_4334_67;
  assign T_23676_39 = T_4334_117;
  assign T_23676_40 = T_4334_147;
  assign T_23676_41 = T_4334_72;
  assign T_23676_42 = T_4334_35;
  assign T_23676_43 = T_4334_146;
  assign T_23676_44 = T_4334_112;
  assign T_23676_45 = T_4334_76;
  assign T_23676_46 = T_4334_61;
  assign T_23676_47 = T_4334_156;
  assign T_23676_48 = T_4334_120;
  assign T_23676_49 = T_4334_115;
  assign T_23676_50 = T_4334_142;
  assign T_23676_51 = T_4334_153;
  assign T_23676_52 = 1'h1;
  assign T_23676_53 = 1'h1;
  assign T_23676_54 = 1'h1;
  assign T_23676_55 = 1'h1;
  assign T_23676_56 = 1'h1;
  assign T_23676_57 = 1'h1;
  assign T_23676_58 = 1'h1;
  assign T_23676_59 = 1'h1;
  assign T_23676_60 = 1'h1;
  assign T_23676_61 = 1'h1;
  assign T_23676_62 = 1'h1;
  assign T_23676_63 = 1'h1;
  assign T_23676_64 = T_21743;
  assign T_23676_65 = T_21766;
  assign T_23676_66 = 1'h1;
  assign T_23676_67 = 1'h1;
  assign T_23676_68 = 1'h1;
  assign T_23676_69 = 1'h1;
  assign T_23676_70 = 1'h1;
  assign T_23676_71 = 1'h1;
  assign T_23676_72 = 1'h1;
  assign T_23676_73 = 1'h1;
  assign T_23676_74 = 1'h1;
  assign T_23676_75 = 1'h1;
  assign T_23676_76 = 1'h1;
  assign T_23676_77 = 1'h1;
  assign T_23676_78 = 1'h1;
  assign T_23676_79 = 1'h1;
  assign T_23676_80 = 1'h1;
  assign T_23676_81 = 1'h1;
  assign T_23676_82 = 1'h1;
  assign T_23676_83 = 1'h1;
  assign T_23676_84 = 1'h1;
  assign T_23676_85 = 1'h1;
  assign T_23676_86 = 1'h1;
  assign T_23676_87 = 1'h1;
  assign T_23676_88 = 1'h1;
  assign T_23676_89 = 1'h1;
  assign T_23676_90 = 1'h1;
  assign T_23676_91 = 1'h1;
  assign T_23676_92 = 1'h1;
  assign T_23676_93 = 1'h1;
  assign T_23676_94 = 1'h1;
  assign T_23676_95 = 1'h1;
  assign T_23676_96 = 1'h1;
  assign T_23676_97 = 1'h1;
  assign T_23676_98 = 1'h1;
  assign T_23676_99 = 1'h1;
  assign T_23676_100 = 1'h1;
  assign T_23676_101 = 1'h1;
  assign T_23676_102 = 1'h1;
  assign T_23676_103 = 1'h1;
  assign T_23676_104 = 1'h1;
  assign T_23676_105 = 1'h1;
  assign T_23676_106 = 1'h1;
  assign T_23676_107 = 1'h1;
  assign T_23676_108 = 1'h1;
  assign T_23676_109 = 1'h1;
  assign T_23676_110 = 1'h1;
  assign T_23676_111 = 1'h1;
  assign T_23676_112 = 1'h1;
  assign T_23676_113 = 1'h1;
  assign T_23676_114 = 1'h1;
  assign T_23676_115 = 1'h1;
  assign T_23676_116 = 1'h1;
  assign T_23676_117 = 1'h1;
  assign T_23676_118 = 1'h1;
  assign T_23676_119 = 1'h1;
  assign T_23676_120 = 1'h1;
  assign T_23676_121 = 1'h1;
  assign T_23676_122 = 1'h1;
  assign T_23676_123 = 1'h1;
  assign T_23676_124 = 1'h1;
  assign T_23676_125 = 1'h1;
  assign T_23676_126 = 1'h1;
  assign T_23676_127 = 1'h1;
  assign T_23676_128 = T_21987;
  assign T_23676_129 = T_22010;
  assign T_23676_130 = 1'h1;
  assign T_23676_131 = 1'h1;
  assign T_23676_132 = 1'h1;
  assign T_23676_133 = 1'h1;
  assign T_23676_134 = 1'h1;
  assign T_23676_135 = 1'h1;
  assign T_23676_136 = 1'h1;
  assign T_23676_137 = 1'h1;
  assign T_23676_138 = 1'h1;
  assign T_23676_139 = 1'h1;
  assign T_23676_140 = 1'h1;
  assign T_23676_141 = 1'h1;
  assign T_23676_142 = 1'h1;
  assign T_23676_143 = 1'h1;
  assign T_23676_144 = 1'h1;
  assign T_23676_145 = 1'h1;
  assign T_23676_146 = 1'h1;
  assign T_23676_147 = 1'h1;
  assign T_23676_148 = 1'h1;
  assign T_23676_149 = 1'h1;
  assign T_23676_150 = 1'h1;
  assign T_23676_151 = 1'h1;
  assign T_23676_152 = 1'h1;
  assign T_23676_153 = 1'h1;
  assign T_23676_154 = 1'h1;
  assign T_23676_155 = 1'h1;
  assign T_23676_156 = 1'h1;
  assign T_23676_157 = 1'h1;
  assign T_23676_158 = 1'h1;
  assign T_23676_159 = 1'h1;
  assign T_23676_160 = 1'h1;
  assign T_23676_161 = 1'h1;
  assign T_23676_162 = 1'h1;
  assign T_23676_163 = 1'h1;
  assign T_23676_164 = 1'h1;
  assign T_23676_165 = 1'h1;
  assign T_23676_166 = 1'h1;
  assign T_23676_167 = 1'h1;
  assign T_23676_168 = 1'h1;
  assign T_23676_169 = 1'h1;
  assign T_23676_170 = 1'h1;
  assign T_23676_171 = 1'h1;
  assign T_23676_172 = 1'h1;
  assign T_23676_173 = 1'h1;
  assign T_23676_174 = 1'h1;
  assign T_23676_175 = 1'h1;
  assign T_23676_176 = 1'h1;
  assign T_23676_177 = 1'h1;
  assign T_23676_178 = 1'h1;
  assign T_23676_179 = 1'h1;
  assign T_23676_180 = 1'h1;
  assign T_23676_181 = 1'h1;
  assign T_23676_182 = 1'h1;
  assign T_23676_183 = 1'h1;
  assign T_23676_184 = 1'h1;
  assign T_23676_185 = 1'h1;
  assign T_23676_186 = 1'h1;
  assign T_23676_187 = 1'h1;
  assign T_23676_188 = 1'h1;
  assign T_23676_189 = 1'h1;
  assign T_23676_190 = 1'h1;
  assign T_23676_191 = 1'h1;
  assign T_23676_192 = 1'h1;
  assign T_23676_193 = 1'h1;
  assign T_23676_194 = 1'h1;
  assign T_23676_195 = 1'h1;
  assign T_23676_196 = 1'h1;
  assign T_23676_197 = 1'h1;
  assign T_23676_198 = 1'h1;
  assign T_23676_199 = 1'h1;
  assign T_23676_200 = 1'h1;
  assign T_23676_201 = 1'h1;
  assign T_23676_202 = 1'h1;
  assign T_23676_203 = 1'h1;
  assign T_23676_204 = 1'h1;
  assign T_23676_205 = 1'h1;
  assign T_23676_206 = 1'h1;
  assign T_23676_207 = 1'h1;
  assign T_23676_208 = 1'h1;
  assign T_23676_209 = 1'h1;
  assign T_23676_210 = 1'h1;
  assign T_23676_211 = 1'h1;
  assign T_23676_212 = 1'h1;
  assign T_23676_213 = 1'h1;
  assign T_23676_214 = 1'h1;
  assign T_23676_215 = 1'h1;
  assign T_23676_216 = 1'h1;
  assign T_23676_217 = 1'h1;
  assign T_23676_218 = 1'h1;
  assign T_23676_219 = 1'h1;
  assign T_23676_220 = 1'h1;
  assign T_23676_221 = 1'h1;
  assign T_23676_222 = 1'h1;
  assign T_23676_223 = 1'h1;
  assign T_23676_224 = 1'h1;
  assign T_23676_225 = 1'h1;
  assign T_23676_226 = 1'h1;
  assign T_23676_227 = 1'h1;
  assign T_23676_228 = 1'h1;
  assign T_23676_229 = 1'h1;
  assign T_23676_230 = 1'h1;
  assign T_23676_231 = 1'h1;
  assign T_23676_232 = 1'h1;
  assign T_23676_233 = 1'h1;
  assign T_23676_234 = 1'h1;
  assign T_23676_235 = 1'h1;
  assign T_23676_236 = 1'h1;
  assign T_23676_237 = 1'h1;
  assign T_23676_238 = 1'h1;
  assign T_23676_239 = 1'h1;
  assign T_23676_240 = 1'h1;
  assign T_23676_241 = 1'h1;
  assign T_23676_242 = 1'h1;
  assign T_23676_243 = 1'h1;
  assign T_23676_244 = 1'h1;
  assign T_23676_245 = 1'h1;
  assign T_23676_246 = 1'h1;
  assign T_23676_247 = 1'h1;
  assign T_23676_248 = 1'h1;
  assign T_23676_249 = 1'h1;
  assign T_23676_250 = 1'h1;
  assign T_23676_251 = 1'h1;
  assign T_23676_252 = 1'h1;
  assign T_23676_253 = 1'h1;
  assign T_23676_254 = 1'h1;
  assign T_23676_255 = 1'h1;
  assign T_23676_256 = T_4334_78;
  assign T_23676_257 = T_4334_63;
  assign T_23676_258 = 1'h1;
  assign T_23676_259 = 1'h1;
  assign T_23676_260 = 1'h1;
  assign T_23676_261 = 1'h1;
  assign T_23676_262 = 1'h1;
  assign T_23676_263 = 1'h1;
  assign T_23676_264 = 1'h1;
  assign T_23676_265 = 1'h1;
  assign T_23676_266 = 1'h1;
  assign T_23676_267 = 1'h1;
  assign T_23676_268 = 1'h1;
  assign T_23676_269 = 1'h1;
  assign T_23676_270 = 1'h1;
  assign T_23676_271 = 1'h1;
  assign T_23676_272 = 1'h1;
  assign T_23676_273 = 1'h1;
  assign T_23676_274 = 1'h1;
  assign T_23676_275 = 1'h1;
  assign T_23676_276 = 1'h1;
  assign T_23676_277 = 1'h1;
  assign T_23676_278 = 1'h1;
  assign T_23676_279 = 1'h1;
  assign T_23676_280 = 1'h1;
  assign T_23676_281 = 1'h1;
  assign T_23676_282 = 1'h1;
  assign T_23676_283 = 1'h1;
  assign T_23676_284 = 1'h1;
  assign T_23676_285 = 1'h1;
  assign T_23676_286 = 1'h1;
  assign T_23676_287 = 1'h1;
  assign T_23676_288 = 1'h1;
  assign T_23676_289 = 1'h1;
  assign T_23676_290 = 1'h1;
  assign T_23676_291 = 1'h1;
  assign T_23676_292 = 1'h1;
  assign T_23676_293 = 1'h1;
  assign T_23676_294 = 1'h1;
  assign T_23676_295 = 1'h1;
  assign T_23676_296 = 1'h1;
  assign T_23676_297 = 1'h1;
  assign T_23676_298 = 1'h1;
  assign T_23676_299 = 1'h1;
  assign T_23676_300 = 1'h1;
  assign T_23676_301 = 1'h1;
  assign T_23676_302 = 1'h1;
  assign T_23676_303 = 1'h1;
  assign T_23676_304 = 1'h1;
  assign T_23676_305 = 1'h1;
  assign T_23676_306 = 1'h1;
  assign T_23676_307 = 1'h1;
  assign T_23676_308 = 1'h1;
  assign T_23676_309 = 1'h1;
  assign T_23676_310 = 1'h1;
  assign T_23676_311 = 1'h1;
  assign T_23676_312 = 1'h1;
  assign T_23676_313 = 1'h1;
  assign T_23676_314 = 1'h1;
  assign T_23676_315 = 1'h1;
  assign T_23676_316 = 1'h1;
  assign T_23676_317 = 1'h1;
  assign T_23676_318 = 1'h1;
  assign T_23676_319 = 1'h1;
  assign T_23676_320 = 1'h1;
  assign T_23676_321 = 1'h1;
  assign T_23676_322 = 1'h1;
  assign T_23676_323 = 1'h1;
  assign T_23676_324 = 1'h1;
  assign T_23676_325 = 1'h1;
  assign T_23676_326 = 1'h1;
  assign T_23676_327 = 1'h1;
  assign T_23676_328 = 1'h1;
  assign T_23676_329 = 1'h1;
  assign T_23676_330 = 1'h1;
  assign T_23676_331 = 1'h1;
  assign T_23676_332 = 1'h1;
  assign T_23676_333 = 1'h1;
  assign T_23676_334 = 1'h1;
  assign T_23676_335 = 1'h1;
  assign T_23676_336 = 1'h1;
  assign T_23676_337 = 1'h1;
  assign T_23676_338 = 1'h1;
  assign T_23676_339 = 1'h1;
  assign T_23676_340 = 1'h1;
  assign T_23676_341 = 1'h1;
  assign T_23676_342 = 1'h1;
  assign T_23676_343 = 1'h1;
  assign T_23676_344 = 1'h1;
  assign T_23676_345 = 1'h1;
  assign T_23676_346 = 1'h1;
  assign T_23676_347 = 1'h1;
  assign T_23676_348 = 1'h1;
  assign T_23676_349 = 1'h1;
  assign T_23676_350 = 1'h1;
  assign T_23676_351 = 1'h1;
  assign T_23676_352 = 1'h1;
  assign T_23676_353 = 1'h1;
  assign T_23676_354 = 1'h1;
  assign T_23676_355 = 1'h1;
  assign T_23676_356 = 1'h1;
  assign T_23676_357 = 1'h1;
  assign T_23676_358 = 1'h1;
  assign T_23676_359 = 1'h1;
  assign T_23676_360 = 1'h1;
  assign T_23676_361 = 1'h1;
  assign T_23676_362 = 1'h1;
  assign T_23676_363 = 1'h1;
  assign T_23676_364 = 1'h1;
  assign T_23676_365 = 1'h1;
  assign T_23676_366 = 1'h1;
  assign T_23676_367 = 1'h1;
  assign T_23676_368 = 1'h1;
  assign T_23676_369 = 1'h1;
  assign T_23676_370 = 1'h1;
  assign T_23676_371 = 1'h1;
  assign T_23676_372 = 1'h1;
  assign T_23676_373 = 1'h1;
  assign T_23676_374 = 1'h1;
  assign T_23676_375 = 1'h1;
  assign T_23676_376 = 1'h1;
  assign T_23676_377 = 1'h1;
  assign T_23676_378 = 1'h1;
  assign T_23676_379 = 1'h1;
  assign T_23676_380 = 1'h1;
  assign T_23676_381 = 1'h1;
  assign T_23676_382 = 1'h1;
  assign T_23676_383 = 1'h1;
  assign T_23676_384 = 1'h1;
  assign T_23676_385 = 1'h1;
  assign T_23676_386 = 1'h1;
  assign T_23676_387 = 1'h1;
  assign T_23676_388 = 1'h1;
  assign T_23676_389 = 1'h1;
  assign T_23676_390 = 1'h1;
  assign T_23676_391 = 1'h1;
  assign T_23676_392 = 1'h1;
  assign T_23676_393 = 1'h1;
  assign T_23676_394 = 1'h1;
  assign T_23676_395 = 1'h1;
  assign T_23676_396 = 1'h1;
  assign T_23676_397 = 1'h1;
  assign T_23676_398 = 1'h1;
  assign T_23676_399 = 1'h1;
  assign T_23676_400 = 1'h1;
  assign T_23676_401 = 1'h1;
  assign T_23676_402 = 1'h1;
  assign T_23676_403 = 1'h1;
  assign T_23676_404 = 1'h1;
  assign T_23676_405 = 1'h1;
  assign T_23676_406 = 1'h1;
  assign T_23676_407 = 1'h1;
  assign T_23676_408 = 1'h1;
  assign T_23676_409 = 1'h1;
  assign T_23676_410 = 1'h1;
  assign T_23676_411 = 1'h1;
  assign T_23676_412 = 1'h1;
  assign T_23676_413 = 1'h1;
  assign T_23676_414 = 1'h1;
  assign T_23676_415 = 1'h1;
  assign T_23676_416 = 1'h1;
  assign T_23676_417 = 1'h1;
  assign T_23676_418 = 1'h1;
  assign T_23676_419 = 1'h1;
  assign T_23676_420 = 1'h1;
  assign T_23676_421 = 1'h1;
  assign T_23676_422 = 1'h1;
  assign T_23676_423 = 1'h1;
  assign T_23676_424 = 1'h1;
  assign T_23676_425 = 1'h1;
  assign T_23676_426 = 1'h1;
  assign T_23676_427 = 1'h1;
  assign T_23676_428 = 1'h1;
  assign T_23676_429 = 1'h1;
  assign T_23676_430 = 1'h1;
  assign T_23676_431 = 1'h1;
  assign T_23676_432 = 1'h1;
  assign T_23676_433 = 1'h1;
  assign T_23676_434 = 1'h1;
  assign T_23676_435 = 1'h1;
  assign T_23676_436 = 1'h1;
  assign T_23676_437 = 1'h1;
  assign T_23676_438 = 1'h1;
  assign T_23676_439 = 1'h1;
  assign T_23676_440 = 1'h1;
  assign T_23676_441 = 1'h1;
  assign T_23676_442 = 1'h1;
  assign T_23676_443 = 1'h1;
  assign T_23676_444 = 1'h1;
  assign T_23676_445 = 1'h1;
  assign T_23676_446 = 1'h1;
  assign T_23676_447 = 1'h1;
  assign T_23676_448 = 1'h1;
  assign T_23676_449 = 1'h1;
  assign T_23676_450 = 1'h1;
  assign T_23676_451 = 1'h1;
  assign T_23676_452 = 1'h1;
  assign T_23676_453 = 1'h1;
  assign T_23676_454 = 1'h1;
  assign T_23676_455 = 1'h1;
  assign T_23676_456 = 1'h1;
  assign T_23676_457 = 1'h1;
  assign T_23676_458 = 1'h1;
  assign T_23676_459 = 1'h1;
  assign T_23676_460 = 1'h1;
  assign T_23676_461 = 1'h1;
  assign T_23676_462 = 1'h1;
  assign T_23676_463 = 1'h1;
  assign T_23676_464 = 1'h1;
  assign T_23676_465 = 1'h1;
  assign T_23676_466 = 1'h1;
  assign T_23676_467 = 1'h1;
  assign T_23676_468 = 1'h1;
  assign T_23676_469 = 1'h1;
  assign T_23676_470 = 1'h1;
  assign T_23676_471 = 1'h1;
  assign T_23676_472 = 1'h1;
  assign T_23676_473 = 1'h1;
  assign T_23676_474 = 1'h1;
  assign T_23676_475 = 1'h1;
  assign T_23676_476 = 1'h1;
  assign T_23676_477 = 1'h1;
  assign T_23676_478 = 1'h1;
  assign T_23676_479 = 1'h1;
  assign T_23676_480 = 1'h1;
  assign T_23676_481 = 1'h1;
  assign T_23676_482 = 1'h1;
  assign T_23676_483 = 1'h1;
  assign T_23676_484 = 1'h1;
  assign T_23676_485 = 1'h1;
  assign T_23676_486 = 1'h1;
  assign T_23676_487 = 1'h1;
  assign T_23676_488 = 1'h1;
  assign T_23676_489 = 1'h1;
  assign T_23676_490 = 1'h1;
  assign T_23676_491 = 1'h1;
  assign T_23676_492 = 1'h1;
  assign T_23676_493 = 1'h1;
  assign T_23676_494 = 1'h1;
  assign T_23676_495 = 1'h1;
  assign T_23676_496 = 1'h1;
  assign T_23676_497 = 1'h1;
  assign T_23676_498 = 1'h1;
  assign T_23676_499 = 1'h1;
  assign T_23676_500 = 1'h1;
  assign T_23676_501 = 1'h1;
  assign T_23676_502 = 1'h1;
  assign T_23676_503 = 1'h1;
  assign T_23676_504 = 1'h1;
  assign T_23676_505 = 1'h1;
  assign T_23676_506 = 1'h1;
  assign T_23676_507 = 1'h1;
  assign T_23676_508 = 1'h1;
  assign T_23676_509 = 1'h1;
  assign T_23676_510 = 1'h1;
  assign T_23676_511 = 1'h1;
  assign T_24191 = T_3205_bits_index[0];
  assign T_24192 = T_3205_bits_index[1];
  assign T_24193 = T_3205_bits_index[2];
  assign T_24194 = T_3205_bits_index[3];
  assign T_24195 = T_3205_bits_index[4];
  assign T_24196 = T_3205_bits_index[5];
  assign T_24201 = T_3205_bits_index[10];
  assign T_24202 = T_3205_bits_index[11];
  assign T_24210 = T_3205_bits_index[19];
  assign T_24215 = {T_24192,T_24191};
  assign T_24216 = {T_24194,T_24193};
  assign T_24217 = {T_24216,T_24215};
  assign T_24218 = {T_24196,T_24195};
  assign T_24219 = {T_24210,T_24202};
  assign T_24220 = {T_24219,T_24201};
  assign T_24221 = {T_24220,T_24218};
  assign T_24222 = {T_24221,T_24217};
  assign GEN_3 = GEN_933;
  assign GEN_423 = 9'h1 == T_24222 ? T_15504_1 : T_15504_0;
  assign GEN_424 = 9'h2 == T_24222 ? T_15504_2 : GEN_423;
  assign GEN_425 = 9'h3 == T_24222 ? T_15504_3 : GEN_424;
  assign GEN_426 = 9'h4 == T_24222 ? T_15504_4 : GEN_425;
  assign GEN_427 = 9'h5 == T_24222 ? T_15504_5 : GEN_426;
  assign GEN_428 = 9'h6 == T_24222 ? T_15504_6 : GEN_427;
  assign GEN_429 = 9'h7 == T_24222 ? T_15504_7 : GEN_428;
  assign GEN_430 = 9'h8 == T_24222 ? T_15504_8 : GEN_429;
  assign GEN_431 = 9'h9 == T_24222 ? T_15504_9 : GEN_430;
  assign GEN_432 = 9'ha == T_24222 ? T_15504_10 : GEN_431;
  assign GEN_433 = 9'hb == T_24222 ? T_15504_11 : GEN_432;
  assign GEN_434 = 9'hc == T_24222 ? T_15504_12 : GEN_433;
  assign GEN_435 = 9'hd == T_24222 ? T_15504_13 : GEN_434;
  assign GEN_436 = 9'he == T_24222 ? T_15504_14 : GEN_435;
  assign GEN_437 = 9'hf == T_24222 ? T_15504_15 : GEN_436;
  assign GEN_438 = 9'h10 == T_24222 ? T_15504_16 : GEN_437;
  assign GEN_439 = 9'h11 == T_24222 ? T_15504_17 : GEN_438;
  assign GEN_440 = 9'h12 == T_24222 ? T_15504_18 : GEN_439;
  assign GEN_441 = 9'h13 == T_24222 ? T_15504_19 : GEN_440;
  assign GEN_442 = 9'h14 == T_24222 ? T_15504_20 : GEN_441;
  assign GEN_443 = 9'h15 == T_24222 ? T_15504_21 : GEN_442;
  assign GEN_444 = 9'h16 == T_24222 ? T_15504_22 : GEN_443;
  assign GEN_445 = 9'h17 == T_24222 ? T_15504_23 : GEN_444;
  assign GEN_446 = 9'h18 == T_24222 ? T_15504_24 : GEN_445;
  assign GEN_447 = 9'h19 == T_24222 ? T_15504_25 : GEN_446;
  assign GEN_448 = 9'h1a == T_24222 ? T_15504_26 : GEN_447;
  assign GEN_449 = 9'h1b == T_24222 ? T_15504_27 : GEN_448;
  assign GEN_450 = 9'h1c == T_24222 ? T_15504_28 : GEN_449;
  assign GEN_451 = 9'h1d == T_24222 ? T_15504_29 : GEN_450;
  assign GEN_452 = 9'h1e == T_24222 ? T_15504_30 : GEN_451;
  assign GEN_453 = 9'h1f == T_24222 ? T_15504_31 : GEN_452;
  assign GEN_454 = 9'h20 == T_24222 ? T_15504_32 : GEN_453;
  assign GEN_455 = 9'h21 == T_24222 ? T_15504_33 : GEN_454;
  assign GEN_456 = 9'h22 == T_24222 ? T_15504_34 : GEN_455;
  assign GEN_457 = 9'h23 == T_24222 ? T_15504_35 : GEN_456;
  assign GEN_458 = 9'h24 == T_24222 ? T_15504_36 : GEN_457;
  assign GEN_459 = 9'h25 == T_24222 ? T_15504_37 : GEN_458;
  assign GEN_460 = 9'h26 == T_24222 ? T_15504_38 : GEN_459;
  assign GEN_461 = 9'h27 == T_24222 ? T_15504_39 : GEN_460;
  assign GEN_462 = 9'h28 == T_24222 ? T_15504_40 : GEN_461;
  assign GEN_463 = 9'h29 == T_24222 ? T_15504_41 : GEN_462;
  assign GEN_464 = 9'h2a == T_24222 ? T_15504_42 : GEN_463;
  assign GEN_465 = 9'h2b == T_24222 ? T_15504_43 : GEN_464;
  assign GEN_466 = 9'h2c == T_24222 ? T_15504_44 : GEN_465;
  assign GEN_467 = 9'h2d == T_24222 ? T_15504_45 : GEN_466;
  assign GEN_468 = 9'h2e == T_24222 ? T_15504_46 : GEN_467;
  assign GEN_469 = 9'h2f == T_24222 ? T_15504_47 : GEN_468;
  assign GEN_470 = 9'h30 == T_24222 ? T_15504_48 : GEN_469;
  assign GEN_471 = 9'h31 == T_24222 ? T_15504_49 : GEN_470;
  assign GEN_472 = 9'h32 == T_24222 ? T_15504_50 : GEN_471;
  assign GEN_473 = 9'h33 == T_24222 ? T_15504_51 : GEN_472;
  assign GEN_474 = 9'h34 == T_24222 ? T_15504_52 : GEN_473;
  assign GEN_475 = 9'h35 == T_24222 ? T_15504_53 : GEN_474;
  assign GEN_476 = 9'h36 == T_24222 ? T_15504_54 : GEN_475;
  assign GEN_477 = 9'h37 == T_24222 ? T_15504_55 : GEN_476;
  assign GEN_478 = 9'h38 == T_24222 ? T_15504_56 : GEN_477;
  assign GEN_479 = 9'h39 == T_24222 ? T_15504_57 : GEN_478;
  assign GEN_480 = 9'h3a == T_24222 ? T_15504_58 : GEN_479;
  assign GEN_481 = 9'h3b == T_24222 ? T_15504_59 : GEN_480;
  assign GEN_482 = 9'h3c == T_24222 ? T_15504_60 : GEN_481;
  assign GEN_483 = 9'h3d == T_24222 ? T_15504_61 : GEN_482;
  assign GEN_484 = 9'h3e == T_24222 ? T_15504_62 : GEN_483;
  assign GEN_485 = 9'h3f == T_24222 ? T_15504_63 : GEN_484;
  assign GEN_486 = 9'h40 == T_24222 ? T_15504_64 : GEN_485;
  assign GEN_487 = 9'h41 == T_24222 ? T_15504_65 : GEN_486;
  assign GEN_488 = 9'h42 == T_24222 ? T_15504_66 : GEN_487;
  assign GEN_489 = 9'h43 == T_24222 ? T_15504_67 : GEN_488;
  assign GEN_490 = 9'h44 == T_24222 ? T_15504_68 : GEN_489;
  assign GEN_491 = 9'h45 == T_24222 ? T_15504_69 : GEN_490;
  assign GEN_492 = 9'h46 == T_24222 ? T_15504_70 : GEN_491;
  assign GEN_493 = 9'h47 == T_24222 ? T_15504_71 : GEN_492;
  assign GEN_494 = 9'h48 == T_24222 ? T_15504_72 : GEN_493;
  assign GEN_495 = 9'h49 == T_24222 ? T_15504_73 : GEN_494;
  assign GEN_496 = 9'h4a == T_24222 ? T_15504_74 : GEN_495;
  assign GEN_497 = 9'h4b == T_24222 ? T_15504_75 : GEN_496;
  assign GEN_498 = 9'h4c == T_24222 ? T_15504_76 : GEN_497;
  assign GEN_499 = 9'h4d == T_24222 ? T_15504_77 : GEN_498;
  assign GEN_500 = 9'h4e == T_24222 ? T_15504_78 : GEN_499;
  assign GEN_501 = 9'h4f == T_24222 ? T_15504_79 : GEN_500;
  assign GEN_502 = 9'h50 == T_24222 ? T_15504_80 : GEN_501;
  assign GEN_503 = 9'h51 == T_24222 ? T_15504_81 : GEN_502;
  assign GEN_504 = 9'h52 == T_24222 ? T_15504_82 : GEN_503;
  assign GEN_505 = 9'h53 == T_24222 ? T_15504_83 : GEN_504;
  assign GEN_506 = 9'h54 == T_24222 ? T_15504_84 : GEN_505;
  assign GEN_507 = 9'h55 == T_24222 ? T_15504_85 : GEN_506;
  assign GEN_508 = 9'h56 == T_24222 ? T_15504_86 : GEN_507;
  assign GEN_509 = 9'h57 == T_24222 ? T_15504_87 : GEN_508;
  assign GEN_510 = 9'h58 == T_24222 ? T_15504_88 : GEN_509;
  assign GEN_511 = 9'h59 == T_24222 ? T_15504_89 : GEN_510;
  assign GEN_512 = 9'h5a == T_24222 ? T_15504_90 : GEN_511;
  assign GEN_513 = 9'h5b == T_24222 ? T_15504_91 : GEN_512;
  assign GEN_514 = 9'h5c == T_24222 ? T_15504_92 : GEN_513;
  assign GEN_515 = 9'h5d == T_24222 ? T_15504_93 : GEN_514;
  assign GEN_516 = 9'h5e == T_24222 ? T_15504_94 : GEN_515;
  assign GEN_517 = 9'h5f == T_24222 ? T_15504_95 : GEN_516;
  assign GEN_518 = 9'h60 == T_24222 ? T_15504_96 : GEN_517;
  assign GEN_519 = 9'h61 == T_24222 ? T_15504_97 : GEN_518;
  assign GEN_520 = 9'h62 == T_24222 ? T_15504_98 : GEN_519;
  assign GEN_521 = 9'h63 == T_24222 ? T_15504_99 : GEN_520;
  assign GEN_522 = 9'h64 == T_24222 ? T_15504_100 : GEN_521;
  assign GEN_523 = 9'h65 == T_24222 ? T_15504_101 : GEN_522;
  assign GEN_524 = 9'h66 == T_24222 ? T_15504_102 : GEN_523;
  assign GEN_525 = 9'h67 == T_24222 ? T_15504_103 : GEN_524;
  assign GEN_526 = 9'h68 == T_24222 ? T_15504_104 : GEN_525;
  assign GEN_527 = 9'h69 == T_24222 ? T_15504_105 : GEN_526;
  assign GEN_528 = 9'h6a == T_24222 ? T_15504_106 : GEN_527;
  assign GEN_529 = 9'h6b == T_24222 ? T_15504_107 : GEN_528;
  assign GEN_530 = 9'h6c == T_24222 ? T_15504_108 : GEN_529;
  assign GEN_531 = 9'h6d == T_24222 ? T_15504_109 : GEN_530;
  assign GEN_532 = 9'h6e == T_24222 ? T_15504_110 : GEN_531;
  assign GEN_533 = 9'h6f == T_24222 ? T_15504_111 : GEN_532;
  assign GEN_534 = 9'h70 == T_24222 ? T_15504_112 : GEN_533;
  assign GEN_535 = 9'h71 == T_24222 ? T_15504_113 : GEN_534;
  assign GEN_536 = 9'h72 == T_24222 ? T_15504_114 : GEN_535;
  assign GEN_537 = 9'h73 == T_24222 ? T_15504_115 : GEN_536;
  assign GEN_538 = 9'h74 == T_24222 ? T_15504_116 : GEN_537;
  assign GEN_539 = 9'h75 == T_24222 ? T_15504_117 : GEN_538;
  assign GEN_540 = 9'h76 == T_24222 ? T_15504_118 : GEN_539;
  assign GEN_541 = 9'h77 == T_24222 ? T_15504_119 : GEN_540;
  assign GEN_542 = 9'h78 == T_24222 ? T_15504_120 : GEN_541;
  assign GEN_543 = 9'h79 == T_24222 ? T_15504_121 : GEN_542;
  assign GEN_544 = 9'h7a == T_24222 ? T_15504_122 : GEN_543;
  assign GEN_545 = 9'h7b == T_24222 ? T_15504_123 : GEN_544;
  assign GEN_546 = 9'h7c == T_24222 ? T_15504_124 : GEN_545;
  assign GEN_547 = 9'h7d == T_24222 ? T_15504_125 : GEN_546;
  assign GEN_548 = 9'h7e == T_24222 ? T_15504_126 : GEN_547;
  assign GEN_549 = 9'h7f == T_24222 ? T_15504_127 : GEN_548;
  assign GEN_550 = 9'h80 == T_24222 ? T_15504_128 : GEN_549;
  assign GEN_551 = 9'h81 == T_24222 ? T_15504_129 : GEN_550;
  assign GEN_552 = 9'h82 == T_24222 ? T_15504_130 : GEN_551;
  assign GEN_553 = 9'h83 == T_24222 ? T_15504_131 : GEN_552;
  assign GEN_554 = 9'h84 == T_24222 ? T_15504_132 : GEN_553;
  assign GEN_555 = 9'h85 == T_24222 ? T_15504_133 : GEN_554;
  assign GEN_556 = 9'h86 == T_24222 ? T_15504_134 : GEN_555;
  assign GEN_557 = 9'h87 == T_24222 ? T_15504_135 : GEN_556;
  assign GEN_558 = 9'h88 == T_24222 ? T_15504_136 : GEN_557;
  assign GEN_559 = 9'h89 == T_24222 ? T_15504_137 : GEN_558;
  assign GEN_560 = 9'h8a == T_24222 ? T_15504_138 : GEN_559;
  assign GEN_561 = 9'h8b == T_24222 ? T_15504_139 : GEN_560;
  assign GEN_562 = 9'h8c == T_24222 ? T_15504_140 : GEN_561;
  assign GEN_563 = 9'h8d == T_24222 ? T_15504_141 : GEN_562;
  assign GEN_564 = 9'h8e == T_24222 ? T_15504_142 : GEN_563;
  assign GEN_565 = 9'h8f == T_24222 ? T_15504_143 : GEN_564;
  assign GEN_566 = 9'h90 == T_24222 ? T_15504_144 : GEN_565;
  assign GEN_567 = 9'h91 == T_24222 ? T_15504_145 : GEN_566;
  assign GEN_568 = 9'h92 == T_24222 ? T_15504_146 : GEN_567;
  assign GEN_569 = 9'h93 == T_24222 ? T_15504_147 : GEN_568;
  assign GEN_570 = 9'h94 == T_24222 ? T_15504_148 : GEN_569;
  assign GEN_571 = 9'h95 == T_24222 ? T_15504_149 : GEN_570;
  assign GEN_572 = 9'h96 == T_24222 ? T_15504_150 : GEN_571;
  assign GEN_573 = 9'h97 == T_24222 ? T_15504_151 : GEN_572;
  assign GEN_574 = 9'h98 == T_24222 ? T_15504_152 : GEN_573;
  assign GEN_575 = 9'h99 == T_24222 ? T_15504_153 : GEN_574;
  assign GEN_576 = 9'h9a == T_24222 ? T_15504_154 : GEN_575;
  assign GEN_577 = 9'h9b == T_24222 ? T_15504_155 : GEN_576;
  assign GEN_578 = 9'h9c == T_24222 ? T_15504_156 : GEN_577;
  assign GEN_579 = 9'h9d == T_24222 ? T_15504_157 : GEN_578;
  assign GEN_580 = 9'h9e == T_24222 ? T_15504_158 : GEN_579;
  assign GEN_581 = 9'h9f == T_24222 ? T_15504_159 : GEN_580;
  assign GEN_582 = 9'ha0 == T_24222 ? T_15504_160 : GEN_581;
  assign GEN_583 = 9'ha1 == T_24222 ? T_15504_161 : GEN_582;
  assign GEN_584 = 9'ha2 == T_24222 ? T_15504_162 : GEN_583;
  assign GEN_585 = 9'ha3 == T_24222 ? T_15504_163 : GEN_584;
  assign GEN_586 = 9'ha4 == T_24222 ? T_15504_164 : GEN_585;
  assign GEN_587 = 9'ha5 == T_24222 ? T_15504_165 : GEN_586;
  assign GEN_588 = 9'ha6 == T_24222 ? T_15504_166 : GEN_587;
  assign GEN_589 = 9'ha7 == T_24222 ? T_15504_167 : GEN_588;
  assign GEN_590 = 9'ha8 == T_24222 ? T_15504_168 : GEN_589;
  assign GEN_591 = 9'ha9 == T_24222 ? T_15504_169 : GEN_590;
  assign GEN_592 = 9'haa == T_24222 ? T_15504_170 : GEN_591;
  assign GEN_593 = 9'hab == T_24222 ? T_15504_171 : GEN_592;
  assign GEN_594 = 9'hac == T_24222 ? T_15504_172 : GEN_593;
  assign GEN_595 = 9'had == T_24222 ? T_15504_173 : GEN_594;
  assign GEN_596 = 9'hae == T_24222 ? T_15504_174 : GEN_595;
  assign GEN_597 = 9'haf == T_24222 ? T_15504_175 : GEN_596;
  assign GEN_598 = 9'hb0 == T_24222 ? T_15504_176 : GEN_597;
  assign GEN_599 = 9'hb1 == T_24222 ? T_15504_177 : GEN_598;
  assign GEN_600 = 9'hb2 == T_24222 ? T_15504_178 : GEN_599;
  assign GEN_601 = 9'hb3 == T_24222 ? T_15504_179 : GEN_600;
  assign GEN_602 = 9'hb4 == T_24222 ? T_15504_180 : GEN_601;
  assign GEN_603 = 9'hb5 == T_24222 ? T_15504_181 : GEN_602;
  assign GEN_604 = 9'hb6 == T_24222 ? T_15504_182 : GEN_603;
  assign GEN_605 = 9'hb7 == T_24222 ? T_15504_183 : GEN_604;
  assign GEN_606 = 9'hb8 == T_24222 ? T_15504_184 : GEN_605;
  assign GEN_607 = 9'hb9 == T_24222 ? T_15504_185 : GEN_606;
  assign GEN_608 = 9'hba == T_24222 ? T_15504_186 : GEN_607;
  assign GEN_609 = 9'hbb == T_24222 ? T_15504_187 : GEN_608;
  assign GEN_610 = 9'hbc == T_24222 ? T_15504_188 : GEN_609;
  assign GEN_611 = 9'hbd == T_24222 ? T_15504_189 : GEN_610;
  assign GEN_612 = 9'hbe == T_24222 ? T_15504_190 : GEN_611;
  assign GEN_613 = 9'hbf == T_24222 ? T_15504_191 : GEN_612;
  assign GEN_614 = 9'hc0 == T_24222 ? T_15504_192 : GEN_613;
  assign GEN_615 = 9'hc1 == T_24222 ? T_15504_193 : GEN_614;
  assign GEN_616 = 9'hc2 == T_24222 ? T_15504_194 : GEN_615;
  assign GEN_617 = 9'hc3 == T_24222 ? T_15504_195 : GEN_616;
  assign GEN_618 = 9'hc4 == T_24222 ? T_15504_196 : GEN_617;
  assign GEN_619 = 9'hc5 == T_24222 ? T_15504_197 : GEN_618;
  assign GEN_620 = 9'hc6 == T_24222 ? T_15504_198 : GEN_619;
  assign GEN_621 = 9'hc7 == T_24222 ? T_15504_199 : GEN_620;
  assign GEN_622 = 9'hc8 == T_24222 ? T_15504_200 : GEN_621;
  assign GEN_623 = 9'hc9 == T_24222 ? T_15504_201 : GEN_622;
  assign GEN_624 = 9'hca == T_24222 ? T_15504_202 : GEN_623;
  assign GEN_625 = 9'hcb == T_24222 ? T_15504_203 : GEN_624;
  assign GEN_626 = 9'hcc == T_24222 ? T_15504_204 : GEN_625;
  assign GEN_627 = 9'hcd == T_24222 ? T_15504_205 : GEN_626;
  assign GEN_628 = 9'hce == T_24222 ? T_15504_206 : GEN_627;
  assign GEN_629 = 9'hcf == T_24222 ? T_15504_207 : GEN_628;
  assign GEN_630 = 9'hd0 == T_24222 ? T_15504_208 : GEN_629;
  assign GEN_631 = 9'hd1 == T_24222 ? T_15504_209 : GEN_630;
  assign GEN_632 = 9'hd2 == T_24222 ? T_15504_210 : GEN_631;
  assign GEN_633 = 9'hd3 == T_24222 ? T_15504_211 : GEN_632;
  assign GEN_634 = 9'hd4 == T_24222 ? T_15504_212 : GEN_633;
  assign GEN_635 = 9'hd5 == T_24222 ? T_15504_213 : GEN_634;
  assign GEN_636 = 9'hd6 == T_24222 ? T_15504_214 : GEN_635;
  assign GEN_637 = 9'hd7 == T_24222 ? T_15504_215 : GEN_636;
  assign GEN_638 = 9'hd8 == T_24222 ? T_15504_216 : GEN_637;
  assign GEN_639 = 9'hd9 == T_24222 ? T_15504_217 : GEN_638;
  assign GEN_640 = 9'hda == T_24222 ? T_15504_218 : GEN_639;
  assign GEN_641 = 9'hdb == T_24222 ? T_15504_219 : GEN_640;
  assign GEN_642 = 9'hdc == T_24222 ? T_15504_220 : GEN_641;
  assign GEN_643 = 9'hdd == T_24222 ? T_15504_221 : GEN_642;
  assign GEN_644 = 9'hde == T_24222 ? T_15504_222 : GEN_643;
  assign GEN_645 = 9'hdf == T_24222 ? T_15504_223 : GEN_644;
  assign GEN_646 = 9'he0 == T_24222 ? T_15504_224 : GEN_645;
  assign GEN_647 = 9'he1 == T_24222 ? T_15504_225 : GEN_646;
  assign GEN_648 = 9'he2 == T_24222 ? T_15504_226 : GEN_647;
  assign GEN_649 = 9'he3 == T_24222 ? T_15504_227 : GEN_648;
  assign GEN_650 = 9'he4 == T_24222 ? T_15504_228 : GEN_649;
  assign GEN_651 = 9'he5 == T_24222 ? T_15504_229 : GEN_650;
  assign GEN_652 = 9'he6 == T_24222 ? T_15504_230 : GEN_651;
  assign GEN_653 = 9'he7 == T_24222 ? T_15504_231 : GEN_652;
  assign GEN_654 = 9'he8 == T_24222 ? T_15504_232 : GEN_653;
  assign GEN_655 = 9'he9 == T_24222 ? T_15504_233 : GEN_654;
  assign GEN_656 = 9'hea == T_24222 ? T_15504_234 : GEN_655;
  assign GEN_657 = 9'heb == T_24222 ? T_15504_235 : GEN_656;
  assign GEN_658 = 9'hec == T_24222 ? T_15504_236 : GEN_657;
  assign GEN_659 = 9'hed == T_24222 ? T_15504_237 : GEN_658;
  assign GEN_660 = 9'hee == T_24222 ? T_15504_238 : GEN_659;
  assign GEN_661 = 9'hef == T_24222 ? T_15504_239 : GEN_660;
  assign GEN_662 = 9'hf0 == T_24222 ? T_15504_240 : GEN_661;
  assign GEN_663 = 9'hf1 == T_24222 ? T_15504_241 : GEN_662;
  assign GEN_664 = 9'hf2 == T_24222 ? T_15504_242 : GEN_663;
  assign GEN_665 = 9'hf3 == T_24222 ? T_15504_243 : GEN_664;
  assign GEN_666 = 9'hf4 == T_24222 ? T_15504_244 : GEN_665;
  assign GEN_667 = 9'hf5 == T_24222 ? T_15504_245 : GEN_666;
  assign GEN_668 = 9'hf6 == T_24222 ? T_15504_246 : GEN_667;
  assign GEN_669 = 9'hf7 == T_24222 ? T_15504_247 : GEN_668;
  assign GEN_670 = 9'hf8 == T_24222 ? T_15504_248 : GEN_669;
  assign GEN_671 = 9'hf9 == T_24222 ? T_15504_249 : GEN_670;
  assign GEN_672 = 9'hfa == T_24222 ? T_15504_250 : GEN_671;
  assign GEN_673 = 9'hfb == T_24222 ? T_15504_251 : GEN_672;
  assign GEN_674 = 9'hfc == T_24222 ? T_15504_252 : GEN_673;
  assign GEN_675 = 9'hfd == T_24222 ? T_15504_253 : GEN_674;
  assign GEN_676 = 9'hfe == T_24222 ? T_15504_254 : GEN_675;
  assign GEN_677 = 9'hff == T_24222 ? T_15504_255 : GEN_676;
  assign GEN_678 = 9'h100 == T_24222 ? T_15504_256 : GEN_677;
  assign GEN_679 = 9'h101 == T_24222 ? T_15504_257 : GEN_678;
  assign GEN_680 = 9'h102 == T_24222 ? T_15504_258 : GEN_679;
  assign GEN_681 = 9'h103 == T_24222 ? T_15504_259 : GEN_680;
  assign GEN_682 = 9'h104 == T_24222 ? T_15504_260 : GEN_681;
  assign GEN_683 = 9'h105 == T_24222 ? T_15504_261 : GEN_682;
  assign GEN_684 = 9'h106 == T_24222 ? T_15504_262 : GEN_683;
  assign GEN_685 = 9'h107 == T_24222 ? T_15504_263 : GEN_684;
  assign GEN_686 = 9'h108 == T_24222 ? T_15504_264 : GEN_685;
  assign GEN_687 = 9'h109 == T_24222 ? T_15504_265 : GEN_686;
  assign GEN_688 = 9'h10a == T_24222 ? T_15504_266 : GEN_687;
  assign GEN_689 = 9'h10b == T_24222 ? T_15504_267 : GEN_688;
  assign GEN_690 = 9'h10c == T_24222 ? T_15504_268 : GEN_689;
  assign GEN_691 = 9'h10d == T_24222 ? T_15504_269 : GEN_690;
  assign GEN_692 = 9'h10e == T_24222 ? T_15504_270 : GEN_691;
  assign GEN_693 = 9'h10f == T_24222 ? T_15504_271 : GEN_692;
  assign GEN_694 = 9'h110 == T_24222 ? T_15504_272 : GEN_693;
  assign GEN_695 = 9'h111 == T_24222 ? T_15504_273 : GEN_694;
  assign GEN_696 = 9'h112 == T_24222 ? T_15504_274 : GEN_695;
  assign GEN_697 = 9'h113 == T_24222 ? T_15504_275 : GEN_696;
  assign GEN_698 = 9'h114 == T_24222 ? T_15504_276 : GEN_697;
  assign GEN_699 = 9'h115 == T_24222 ? T_15504_277 : GEN_698;
  assign GEN_700 = 9'h116 == T_24222 ? T_15504_278 : GEN_699;
  assign GEN_701 = 9'h117 == T_24222 ? T_15504_279 : GEN_700;
  assign GEN_702 = 9'h118 == T_24222 ? T_15504_280 : GEN_701;
  assign GEN_703 = 9'h119 == T_24222 ? T_15504_281 : GEN_702;
  assign GEN_704 = 9'h11a == T_24222 ? T_15504_282 : GEN_703;
  assign GEN_705 = 9'h11b == T_24222 ? T_15504_283 : GEN_704;
  assign GEN_706 = 9'h11c == T_24222 ? T_15504_284 : GEN_705;
  assign GEN_707 = 9'h11d == T_24222 ? T_15504_285 : GEN_706;
  assign GEN_708 = 9'h11e == T_24222 ? T_15504_286 : GEN_707;
  assign GEN_709 = 9'h11f == T_24222 ? T_15504_287 : GEN_708;
  assign GEN_710 = 9'h120 == T_24222 ? T_15504_288 : GEN_709;
  assign GEN_711 = 9'h121 == T_24222 ? T_15504_289 : GEN_710;
  assign GEN_712 = 9'h122 == T_24222 ? T_15504_290 : GEN_711;
  assign GEN_713 = 9'h123 == T_24222 ? T_15504_291 : GEN_712;
  assign GEN_714 = 9'h124 == T_24222 ? T_15504_292 : GEN_713;
  assign GEN_715 = 9'h125 == T_24222 ? T_15504_293 : GEN_714;
  assign GEN_716 = 9'h126 == T_24222 ? T_15504_294 : GEN_715;
  assign GEN_717 = 9'h127 == T_24222 ? T_15504_295 : GEN_716;
  assign GEN_718 = 9'h128 == T_24222 ? T_15504_296 : GEN_717;
  assign GEN_719 = 9'h129 == T_24222 ? T_15504_297 : GEN_718;
  assign GEN_720 = 9'h12a == T_24222 ? T_15504_298 : GEN_719;
  assign GEN_721 = 9'h12b == T_24222 ? T_15504_299 : GEN_720;
  assign GEN_722 = 9'h12c == T_24222 ? T_15504_300 : GEN_721;
  assign GEN_723 = 9'h12d == T_24222 ? T_15504_301 : GEN_722;
  assign GEN_724 = 9'h12e == T_24222 ? T_15504_302 : GEN_723;
  assign GEN_725 = 9'h12f == T_24222 ? T_15504_303 : GEN_724;
  assign GEN_726 = 9'h130 == T_24222 ? T_15504_304 : GEN_725;
  assign GEN_727 = 9'h131 == T_24222 ? T_15504_305 : GEN_726;
  assign GEN_728 = 9'h132 == T_24222 ? T_15504_306 : GEN_727;
  assign GEN_729 = 9'h133 == T_24222 ? T_15504_307 : GEN_728;
  assign GEN_730 = 9'h134 == T_24222 ? T_15504_308 : GEN_729;
  assign GEN_731 = 9'h135 == T_24222 ? T_15504_309 : GEN_730;
  assign GEN_732 = 9'h136 == T_24222 ? T_15504_310 : GEN_731;
  assign GEN_733 = 9'h137 == T_24222 ? T_15504_311 : GEN_732;
  assign GEN_734 = 9'h138 == T_24222 ? T_15504_312 : GEN_733;
  assign GEN_735 = 9'h139 == T_24222 ? T_15504_313 : GEN_734;
  assign GEN_736 = 9'h13a == T_24222 ? T_15504_314 : GEN_735;
  assign GEN_737 = 9'h13b == T_24222 ? T_15504_315 : GEN_736;
  assign GEN_738 = 9'h13c == T_24222 ? T_15504_316 : GEN_737;
  assign GEN_739 = 9'h13d == T_24222 ? T_15504_317 : GEN_738;
  assign GEN_740 = 9'h13e == T_24222 ? T_15504_318 : GEN_739;
  assign GEN_741 = 9'h13f == T_24222 ? T_15504_319 : GEN_740;
  assign GEN_742 = 9'h140 == T_24222 ? T_15504_320 : GEN_741;
  assign GEN_743 = 9'h141 == T_24222 ? T_15504_321 : GEN_742;
  assign GEN_744 = 9'h142 == T_24222 ? T_15504_322 : GEN_743;
  assign GEN_745 = 9'h143 == T_24222 ? T_15504_323 : GEN_744;
  assign GEN_746 = 9'h144 == T_24222 ? T_15504_324 : GEN_745;
  assign GEN_747 = 9'h145 == T_24222 ? T_15504_325 : GEN_746;
  assign GEN_748 = 9'h146 == T_24222 ? T_15504_326 : GEN_747;
  assign GEN_749 = 9'h147 == T_24222 ? T_15504_327 : GEN_748;
  assign GEN_750 = 9'h148 == T_24222 ? T_15504_328 : GEN_749;
  assign GEN_751 = 9'h149 == T_24222 ? T_15504_329 : GEN_750;
  assign GEN_752 = 9'h14a == T_24222 ? T_15504_330 : GEN_751;
  assign GEN_753 = 9'h14b == T_24222 ? T_15504_331 : GEN_752;
  assign GEN_754 = 9'h14c == T_24222 ? T_15504_332 : GEN_753;
  assign GEN_755 = 9'h14d == T_24222 ? T_15504_333 : GEN_754;
  assign GEN_756 = 9'h14e == T_24222 ? T_15504_334 : GEN_755;
  assign GEN_757 = 9'h14f == T_24222 ? T_15504_335 : GEN_756;
  assign GEN_758 = 9'h150 == T_24222 ? T_15504_336 : GEN_757;
  assign GEN_759 = 9'h151 == T_24222 ? T_15504_337 : GEN_758;
  assign GEN_760 = 9'h152 == T_24222 ? T_15504_338 : GEN_759;
  assign GEN_761 = 9'h153 == T_24222 ? T_15504_339 : GEN_760;
  assign GEN_762 = 9'h154 == T_24222 ? T_15504_340 : GEN_761;
  assign GEN_763 = 9'h155 == T_24222 ? T_15504_341 : GEN_762;
  assign GEN_764 = 9'h156 == T_24222 ? T_15504_342 : GEN_763;
  assign GEN_765 = 9'h157 == T_24222 ? T_15504_343 : GEN_764;
  assign GEN_766 = 9'h158 == T_24222 ? T_15504_344 : GEN_765;
  assign GEN_767 = 9'h159 == T_24222 ? T_15504_345 : GEN_766;
  assign GEN_768 = 9'h15a == T_24222 ? T_15504_346 : GEN_767;
  assign GEN_769 = 9'h15b == T_24222 ? T_15504_347 : GEN_768;
  assign GEN_770 = 9'h15c == T_24222 ? T_15504_348 : GEN_769;
  assign GEN_771 = 9'h15d == T_24222 ? T_15504_349 : GEN_770;
  assign GEN_772 = 9'h15e == T_24222 ? T_15504_350 : GEN_771;
  assign GEN_773 = 9'h15f == T_24222 ? T_15504_351 : GEN_772;
  assign GEN_774 = 9'h160 == T_24222 ? T_15504_352 : GEN_773;
  assign GEN_775 = 9'h161 == T_24222 ? T_15504_353 : GEN_774;
  assign GEN_776 = 9'h162 == T_24222 ? T_15504_354 : GEN_775;
  assign GEN_777 = 9'h163 == T_24222 ? T_15504_355 : GEN_776;
  assign GEN_778 = 9'h164 == T_24222 ? T_15504_356 : GEN_777;
  assign GEN_779 = 9'h165 == T_24222 ? T_15504_357 : GEN_778;
  assign GEN_780 = 9'h166 == T_24222 ? T_15504_358 : GEN_779;
  assign GEN_781 = 9'h167 == T_24222 ? T_15504_359 : GEN_780;
  assign GEN_782 = 9'h168 == T_24222 ? T_15504_360 : GEN_781;
  assign GEN_783 = 9'h169 == T_24222 ? T_15504_361 : GEN_782;
  assign GEN_784 = 9'h16a == T_24222 ? T_15504_362 : GEN_783;
  assign GEN_785 = 9'h16b == T_24222 ? T_15504_363 : GEN_784;
  assign GEN_786 = 9'h16c == T_24222 ? T_15504_364 : GEN_785;
  assign GEN_787 = 9'h16d == T_24222 ? T_15504_365 : GEN_786;
  assign GEN_788 = 9'h16e == T_24222 ? T_15504_366 : GEN_787;
  assign GEN_789 = 9'h16f == T_24222 ? T_15504_367 : GEN_788;
  assign GEN_790 = 9'h170 == T_24222 ? T_15504_368 : GEN_789;
  assign GEN_791 = 9'h171 == T_24222 ? T_15504_369 : GEN_790;
  assign GEN_792 = 9'h172 == T_24222 ? T_15504_370 : GEN_791;
  assign GEN_793 = 9'h173 == T_24222 ? T_15504_371 : GEN_792;
  assign GEN_794 = 9'h174 == T_24222 ? T_15504_372 : GEN_793;
  assign GEN_795 = 9'h175 == T_24222 ? T_15504_373 : GEN_794;
  assign GEN_796 = 9'h176 == T_24222 ? T_15504_374 : GEN_795;
  assign GEN_797 = 9'h177 == T_24222 ? T_15504_375 : GEN_796;
  assign GEN_798 = 9'h178 == T_24222 ? T_15504_376 : GEN_797;
  assign GEN_799 = 9'h179 == T_24222 ? T_15504_377 : GEN_798;
  assign GEN_800 = 9'h17a == T_24222 ? T_15504_378 : GEN_799;
  assign GEN_801 = 9'h17b == T_24222 ? T_15504_379 : GEN_800;
  assign GEN_802 = 9'h17c == T_24222 ? T_15504_380 : GEN_801;
  assign GEN_803 = 9'h17d == T_24222 ? T_15504_381 : GEN_802;
  assign GEN_804 = 9'h17e == T_24222 ? T_15504_382 : GEN_803;
  assign GEN_805 = 9'h17f == T_24222 ? T_15504_383 : GEN_804;
  assign GEN_806 = 9'h180 == T_24222 ? T_15504_384 : GEN_805;
  assign GEN_807 = 9'h181 == T_24222 ? T_15504_385 : GEN_806;
  assign GEN_808 = 9'h182 == T_24222 ? T_15504_386 : GEN_807;
  assign GEN_809 = 9'h183 == T_24222 ? T_15504_387 : GEN_808;
  assign GEN_810 = 9'h184 == T_24222 ? T_15504_388 : GEN_809;
  assign GEN_811 = 9'h185 == T_24222 ? T_15504_389 : GEN_810;
  assign GEN_812 = 9'h186 == T_24222 ? T_15504_390 : GEN_811;
  assign GEN_813 = 9'h187 == T_24222 ? T_15504_391 : GEN_812;
  assign GEN_814 = 9'h188 == T_24222 ? T_15504_392 : GEN_813;
  assign GEN_815 = 9'h189 == T_24222 ? T_15504_393 : GEN_814;
  assign GEN_816 = 9'h18a == T_24222 ? T_15504_394 : GEN_815;
  assign GEN_817 = 9'h18b == T_24222 ? T_15504_395 : GEN_816;
  assign GEN_818 = 9'h18c == T_24222 ? T_15504_396 : GEN_817;
  assign GEN_819 = 9'h18d == T_24222 ? T_15504_397 : GEN_818;
  assign GEN_820 = 9'h18e == T_24222 ? T_15504_398 : GEN_819;
  assign GEN_821 = 9'h18f == T_24222 ? T_15504_399 : GEN_820;
  assign GEN_822 = 9'h190 == T_24222 ? T_15504_400 : GEN_821;
  assign GEN_823 = 9'h191 == T_24222 ? T_15504_401 : GEN_822;
  assign GEN_824 = 9'h192 == T_24222 ? T_15504_402 : GEN_823;
  assign GEN_825 = 9'h193 == T_24222 ? T_15504_403 : GEN_824;
  assign GEN_826 = 9'h194 == T_24222 ? T_15504_404 : GEN_825;
  assign GEN_827 = 9'h195 == T_24222 ? T_15504_405 : GEN_826;
  assign GEN_828 = 9'h196 == T_24222 ? T_15504_406 : GEN_827;
  assign GEN_829 = 9'h197 == T_24222 ? T_15504_407 : GEN_828;
  assign GEN_830 = 9'h198 == T_24222 ? T_15504_408 : GEN_829;
  assign GEN_831 = 9'h199 == T_24222 ? T_15504_409 : GEN_830;
  assign GEN_832 = 9'h19a == T_24222 ? T_15504_410 : GEN_831;
  assign GEN_833 = 9'h19b == T_24222 ? T_15504_411 : GEN_832;
  assign GEN_834 = 9'h19c == T_24222 ? T_15504_412 : GEN_833;
  assign GEN_835 = 9'h19d == T_24222 ? T_15504_413 : GEN_834;
  assign GEN_836 = 9'h19e == T_24222 ? T_15504_414 : GEN_835;
  assign GEN_837 = 9'h19f == T_24222 ? T_15504_415 : GEN_836;
  assign GEN_838 = 9'h1a0 == T_24222 ? T_15504_416 : GEN_837;
  assign GEN_839 = 9'h1a1 == T_24222 ? T_15504_417 : GEN_838;
  assign GEN_840 = 9'h1a2 == T_24222 ? T_15504_418 : GEN_839;
  assign GEN_841 = 9'h1a3 == T_24222 ? T_15504_419 : GEN_840;
  assign GEN_842 = 9'h1a4 == T_24222 ? T_15504_420 : GEN_841;
  assign GEN_843 = 9'h1a5 == T_24222 ? T_15504_421 : GEN_842;
  assign GEN_844 = 9'h1a6 == T_24222 ? T_15504_422 : GEN_843;
  assign GEN_845 = 9'h1a7 == T_24222 ? T_15504_423 : GEN_844;
  assign GEN_846 = 9'h1a8 == T_24222 ? T_15504_424 : GEN_845;
  assign GEN_847 = 9'h1a9 == T_24222 ? T_15504_425 : GEN_846;
  assign GEN_848 = 9'h1aa == T_24222 ? T_15504_426 : GEN_847;
  assign GEN_849 = 9'h1ab == T_24222 ? T_15504_427 : GEN_848;
  assign GEN_850 = 9'h1ac == T_24222 ? T_15504_428 : GEN_849;
  assign GEN_851 = 9'h1ad == T_24222 ? T_15504_429 : GEN_850;
  assign GEN_852 = 9'h1ae == T_24222 ? T_15504_430 : GEN_851;
  assign GEN_853 = 9'h1af == T_24222 ? T_15504_431 : GEN_852;
  assign GEN_854 = 9'h1b0 == T_24222 ? T_15504_432 : GEN_853;
  assign GEN_855 = 9'h1b1 == T_24222 ? T_15504_433 : GEN_854;
  assign GEN_856 = 9'h1b2 == T_24222 ? T_15504_434 : GEN_855;
  assign GEN_857 = 9'h1b3 == T_24222 ? T_15504_435 : GEN_856;
  assign GEN_858 = 9'h1b4 == T_24222 ? T_15504_436 : GEN_857;
  assign GEN_859 = 9'h1b5 == T_24222 ? T_15504_437 : GEN_858;
  assign GEN_860 = 9'h1b6 == T_24222 ? T_15504_438 : GEN_859;
  assign GEN_861 = 9'h1b7 == T_24222 ? T_15504_439 : GEN_860;
  assign GEN_862 = 9'h1b8 == T_24222 ? T_15504_440 : GEN_861;
  assign GEN_863 = 9'h1b9 == T_24222 ? T_15504_441 : GEN_862;
  assign GEN_864 = 9'h1ba == T_24222 ? T_15504_442 : GEN_863;
  assign GEN_865 = 9'h1bb == T_24222 ? T_15504_443 : GEN_864;
  assign GEN_866 = 9'h1bc == T_24222 ? T_15504_444 : GEN_865;
  assign GEN_867 = 9'h1bd == T_24222 ? T_15504_445 : GEN_866;
  assign GEN_868 = 9'h1be == T_24222 ? T_15504_446 : GEN_867;
  assign GEN_869 = 9'h1bf == T_24222 ? T_15504_447 : GEN_868;
  assign GEN_870 = 9'h1c0 == T_24222 ? T_15504_448 : GEN_869;
  assign GEN_871 = 9'h1c1 == T_24222 ? T_15504_449 : GEN_870;
  assign GEN_872 = 9'h1c2 == T_24222 ? T_15504_450 : GEN_871;
  assign GEN_873 = 9'h1c3 == T_24222 ? T_15504_451 : GEN_872;
  assign GEN_874 = 9'h1c4 == T_24222 ? T_15504_452 : GEN_873;
  assign GEN_875 = 9'h1c5 == T_24222 ? T_15504_453 : GEN_874;
  assign GEN_876 = 9'h1c6 == T_24222 ? T_15504_454 : GEN_875;
  assign GEN_877 = 9'h1c7 == T_24222 ? T_15504_455 : GEN_876;
  assign GEN_878 = 9'h1c8 == T_24222 ? T_15504_456 : GEN_877;
  assign GEN_879 = 9'h1c9 == T_24222 ? T_15504_457 : GEN_878;
  assign GEN_880 = 9'h1ca == T_24222 ? T_15504_458 : GEN_879;
  assign GEN_881 = 9'h1cb == T_24222 ? T_15504_459 : GEN_880;
  assign GEN_882 = 9'h1cc == T_24222 ? T_15504_460 : GEN_881;
  assign GEN_883 = 9'h1cd == T_24222 ? T_15504_461 : GEN_882;
  assign GEN_884 = 9'h1ce == T_24222 ? T_15504_462 : GEN_883;
  assign GEN_885 = 9'h1cf == T_24222 ? T_15504_463 : GEN_884;
  assign GEN_886 = 9'h1d0 == T_24222 ? T_15504_464 : GEN_885;
  assign GEN_887 = 9'h1d1 == T_24222 ? T_15504_465 : GEN_886;
  assign GEN_888 = 9'h1d2 == T_24222 ? T_15504_466 : GEN_887;
  assign GEN_889 = 9'h1d3 == T_24222 ? T_15504_467 : GEN_888;
  assign GEN_890 = 9'h1d4 == T_24222 ? T_15504_468 : GEN_889;
  assign GEN_891 = 9'h1d5 == T_24222 ? T_15504_469 : GEN_890;
  assign GEN_892 = 9'h1d6 == T_24222 ? T_15504_470 : GEN_891;
  assign GEN_893 = 9'h1d7 == T_24222 ? T_15504_471 : GEN_892;
  assign GEN_894 = 9'h1d8 == T_24222 ? T_15504_472 : GEN_893;
  assign GEN_895 = 9'h1d9 == T_24222 ? T_15504_473 : GEN_894;
  assign GEN_896 = 9'h1da == T_24222 ? T_15504_474 : GEN_895;
  assign GEN_897 = 9'h1db == T_24222 ? T_15504_475 : GEN_896;
  assign GEN_898 = 9'h1dc == T_24222 ? T_15504_476 : GEN_897;
  assign GEN_899 = 9'h1dd == T_24222 ? T_15504_477 : GEN_898;
  assign GEN_900 = 9'h1de == T_24222 ? T_15504_478 : GEN_899;
  assign GEN_901 = 9'h1df == T_24222 ? T_15504_479 : GEN_900;
  assign GEN_902 = 9'h1e0 == T_24222 ? T_15504_480 : GEN_901;
  assign GEN_903 = 9'h1e1 == T_24222 ? T_15504_481 : GEN_902;
  assign GEN_904 = 9'h1e2 == T_24222 ? T_15504_482 : GEN_903;
  assign GEN_905 = 9'h1e3 == T_24222 ? T_15504_483 : GEN_904;
  assign GEN_906 = 9'h1e4 == T_24222 ? T_15504_484 : GEN_905;
  assign GEN_907 = 9'h1e5 == T_24222 ? T_15504_485 : GEN_906;
  assign GEN_908 = 9'h1e6 == T_24222 ? T_15504_486 : GEN_907;
  assign GEN_909 = 9'h1e7 == T_24222 ? T_15504_487 : GEN_908;
  assign GEN_910 = 9'h1e8 == T_24222 ? T_15504_488 : GEN_909;
  assign GEN_911 = 9'h1e9 == T_24222 ? T_15504_489 : GEN_910;
  assign GEN_912 = 9'h1ea == T_24222 ? T_15504_490 : GEN_911;
  assign GEN_913 = 9'h1eb == T_24222 ? T_15504_491 : GEN_912;
  assign GEN_914 = 9'h1ec == T_24222 ? T_15504_492 : GEN_913;
  assign GEN_915 = 9'h1ed == T_24222 ? T_15504_493 : GEN_914;
  assign GEN_916 = 9'h1ee == T_24222 ? T_15504_494 : GEN_915;
  assign GEN_917 = 9'h1ef == T_24222 ? T_15504_495 : GEN_916;
  assign GEN_918 = 9'h1f0 == T_24222 ? T_15504_496 : GEN_917;
  assign GEN_919 = 9'h1f1 == T_24222 ? T_15504_497 : GEN_918;
  assign GEN_920 = 9'h1f2 == T_24222 ? T_15504_498 : GEN_919;
  assign GEN_921 = 9'h1f3 == T_24222 ? T_15504_499 : GEN_920;
  assign GEN_922 = 9'h1f4 == T_24222 ? T_15504_500 : GEN_921;
  assign GEN_923 = 9'h1f5 == T_24222 ? T_15504_501 : GEN_922;
  assign GEN_924 = 9'h1f6 == T_24222 ? T_15504_502 : GEN_923;
  assign GEN_925 = 9'h1f7 == T_24222 ? T_15504_503 : GEN_924;
  assign GEN_926 = 9'h1f8 == T_24222 ? T_15504_504 : GEN_925;
  assign GEN_927 = 9'h1f9 == T_24222 ? T_15504_505 : GEN_926;
  assign GEN_928 = 9'h1fa == T_24222 ? T_15504_506 : GEN_927;
  assign GEN_929 = 9'h1fb == T_24222 ? T_15504_507 : GEN_928;
  assign GEN_930 = 9'h1fc == T_24222 ? T_15504_508 : GEN_929;
  assign GEN_931 = 9'h1fd == T_24222 ? T_15504_509 : GEN_930;
  assign GEN_932 = 9'h1fe == T_24222 ? T_15504_510 : GEN_931;
  assign GEN_933 = 9'h1ff == T_24222 ? T_15504_511 : GEN_932;
  assign GEN_4 = GEN_1444;
  assign GEN_934 = 9'h1 == T_24222 ? T_18228_1 : T_18228_0;
  assign GEN_935 = 9'h2 == T_24222 ? T_18228_2 : GEN_934;
  assign GEN_936 = 9'h3 == T_24222 ? T_18228_3 : GEN_935;
  assign GEN_937 = 9'h4 == T_24222 ? T_18228_4 : GEN_936;
  assign GEN_938 = 9'h5 == T_24222 ? T_18228_5 : GEN_937;
  assign GEN_939 = 9'h6 == T_24222 ? T_18228_6 : GEN_938;
  assign GEN_940 = 9'h7 == T_24222 ? T_18228_7 : GEN_939;
  assign GEN_941 = 9'h8 == T_24222 ? T_18228_8 : GEN_940;
  assign GEN_942 = 9'h9 == T_24222 ? T_18228_9 : GEN_941;
  assign GEN_943 = 9'ha == T_24222 ? T_18228_10 : GEN_942;
  assign GEN_944 = 9'hb == T_24222 ? T_18228_11 : GEN_943;
  assign GEN_945 = 9'hc == T_24222 ? T_18228_12 : GEN_944;
  assign GEN_946 = 9'hd == T_24222 ? T_18228_13 : GEN_945;
  assign GEN_947 = 9'he == T_24222 ? T_18228_14 : GEN_946;
  assign GEN_948 = 9'hf == T_24222 ? T_18228_15 : GEN_947;
  assign GEN_949 = 9'h10 == T_24222 ? T_18228_16 : GEN_948;
  assign GEN_950 = 9'h11 == T_24222 ? T_18228_17 : GEN_949;
  assign GEN_951 = 9'h12 == T_24222 ? T_18228_18 : GEN_950;
  assign GEN_952 = 9'h13 == T_24222 ? T_18228_19 : GEN_951;
  assign GEN_953 = 9'h14 == T_24222 ? T_18228_20 : GEN_952;
  assign GEN_954 = 9'h15 == T_24222 ? T_18228_21 : GEN_953;
  assign GEN_955 = 9'h16 == T_24222 ? T_18228_22 : GEN_954;
  assign GEN_956 = 9'h17 == T_24222 ? T_18228_23 : GEN_955;
  assign GEN_957 = 9'h18 == T_24222 ? T_18228_24 : GEN_956;
  assign GEN_958 = 9'h19 == T_24222 ? T_18228_25 : GEN_957;
  assign GEN_959 = 9'h1a == T_24222 ? T_18228_26 : GEN_958;
  assign GEN_960 = 9'h1b == T_24222 ? T_18228_27 : GEN_959;
  assign GEN_961 = 9'h1c == T_24222 ? T_18228_28 : GEN_960;
  assign GEN_962 = 9'h1d == T_24222 ? T_18228_29 : GEN_961;
  assign GEN_963 = 9'h1e == T_24222 ? T_18228_30 : GEN_962;
  assign GEN_964 = 9'h1f == T_24222 ? T_18228_31 : GEN_963;
  assign GEN_965 = 9'h20 == T_24222 ? T_18228_32 : GEN_964;
  assign GEN_966 = 9'h21 == T_24222 ? T_18228_33 : GEN_965;
  assign GEN_967 = 9'h22 == T_24222 ? T_18228_34 : GEN_966;
  assign GEN_968 = 9'h23 == T_24222 ? T_18228_35 : GEN_967;
  assign GEN_969 = 9'h24 == T_24222 ? T_18228_36 : GEN_968;
  assign GEN_970 = 9'h25 == T_24222 ? T_18228_37 : GEN_969;
  assign GEN_971 = 9'h26 == T_24222 ? T_18228_38 : GEN_970;
  assign GEN_972 = 9'h27 == T_24222 ? T_18228_39 : GEN_971;
  assign GEN_973 = 9'h28 == T_24222 ? T_18228_40 : GEN_972;
  assign GEN_974 = 9'h29 == T_24222 ? T_18228_41 : GEN_973;
  assign GEN_975 = 9'h2a == T_24222 ? T_18228_42 : GEN_974;
  assign GEN_976 = 9'h2b == T_24222 ? T_18228_43 : GEN_975;
  assign GEN_977 = 9'h2c == T_24222 ? T_18228_44 : GEN_976;
  assign GEN_978 = 9'h2d == T_24222 ? T_18228_45 : GEN_977;
  assign GEN_979 = 9'h2e == T_24222 ? T_18228_46 : GEN_978;
  assign GEN_980 = 9'h2f == T_24222 ? T_18228_47 : GEN_979;
  assign GEN_981 = 9'h30 == T_24222 ? T_18228_48 : GEN_980;
  assign GEN_982 = 9'h31 == T_24222 ? T_18228_49 : GEN_981;
  assign GEN_983 = 9'h32 == T_24222 ? T_18228_50 : GEN_982;
  assign GEN_984 = 9'h33 == T_24222 ? T_18228_51 : GEN_983;
  assign GEN_985 = 9'h34 == T_24222 ? T_18228_52 : GEN_984;
  assign GEN_986 = 9'h35 == T_24222 ? T_18228_53 : GEN_985;
  assign GEN_987 = 9'h36 == T_24222 ? T_18228_54 : GEN_986;
  assign GEN_988 = 9'h37 == T_24222 ? T_18228_55 : GEN_987;
  assign GEN_989 = 9'h38 == T_24222 ? T_18228_56 : GEN_988;
  assign GEN_990 = 9'h39 == T_24222 ? T_18228_57 : GEN_989;
  assign GEN_991 = 9'h3a == T_24222 ? T_18228_58 : GEN_990;
  assign GEN_992 = 9'h3b == T_24222 ? T_18228_59 : GEN_991;
  assign GEN_993 = 9'h3c == T_24222 ? T_18228_60 : GEN_992;
  assign GEN_994 = 9'h3d == T_24222 ? T_18228_61 : GEN_993;
  assign GEN_995 = 9'h3e == T_24222 ? T_18228_62 : GEN_994;
  assign GEN_996 = 9'h3f == T_24222 ? T_18228_63 : GEN_995;
  assign GEN_997 = 9'h40 == T_24222 ? T_18228_64 : GEN_996;
  assign GEN_998 = 9'h41 == T_24222 ? T_18228_65 : GEN_997;
  assign GEN_999 = 9'h42 == T_24222 ? T_18228_66 : GEN_998;
  assign GEN_1000 = 9'h43 == T_24222 ? T_18228_67 : GEN_999;
  assign GEN_1001 = 9'h44 == T_24222 ? T_18228_68 : GEN_1000;
  assign GEN_1002 = 9'h45 == T_24222 ? T_18228_69 : GEN_1001;
  assign GEN_1003 = 9'h46 == T_24222 ? T_18228_70 : GEN_1002;
  assign GEN_1004 = 9'h47 == T_24222 ? T_18228_71 : GEN_1003;
  assign GEN_1005 = 9'h48 == T_24222 ? T_18228_72 : GEN_1004;
  assign GEN_1006 = 9'h49 == T_24222 ? T_18228_73 : GEN_1005;
  assign GEN_1007 = 9'h4a == T_24222 ? T_18228_74 : GEN_1006;
  assign GEN_1008 = 9'h4b == T_24222 ? T_18228_75 : GEN_1007;
  assign GEN_1009 = 9'h4c == T_24222 ? T_18228_76 : GEN_1008;
  assign GEN_1010 = 9'h4d == T_24222 ? T_18228_77 : GEN_1009;
  assign GEN_1011 = 9'h4e == T_24222 ? T_18228_78 : GEN_1010;
  assign GEN_1012 = 9'h4f == T_24222 ? T_18228_79 : GEN_1011;
  assign GEN_1013 = 9'h50 == T_24222 ? T_18228_80 : GEN_1012;
  assign GEN_1014 = 9'h51 == T_24222 ? T_18228_81 : GEN_1013;
  assign GEN_1015 = 9'h52 == T_24222 ? T_18228_82 : GEN_1014;
  assign GEN_1016 = 9'h53 == T_24222 ? T_18228_83 : GEN_1015;
  assign GEN_1017 = 9'h54 == T_24222 ? T_18228_84 : GEN_1016;
  assign GEN_1018 = 9'h55 == T_24222 ? T_18228_85 : GEN_1017;
  assign GEN_1019 = 9'h56 == T_24222 ? T_18228_86 : GEN_1018;
  assign GEN_1020 = 9'h57 == T_24222 ? T_18228_87 : GEN_1019;
  assign GEN_1021 = 9'h58 == T_24222 ? T_18228_88 : GEN_1020;
  assign GEN_1022 = 9'h59 == T_24222 ? T_18228_89 : GEN_1021;
  assign GEN_1023 = 9'h5a == T_24222 ? T_18228_90 : GEN_1022;
  assign GEN_1024 = 9'h5b == T_24222 ? T_18228_91 : GEN_1023;
  assign GEN_1025 = 9'h5c == T_24222 ? T_18228_92 : GEN_1024;
  assign GEN_1026 = 9'h5d == T_24222 ? T_18228_93 : GEN_1025;
  assign GEN_1027 = 9'h5e == T_24222 ? T_18228_94 : GEN_1026;
  assign GEN_1028 = 9'h5f == T_24222 ? T_18228_95 : GEN_1027;
  assign GEN_1029 = 9'h60 == T_24222 ? T_18228_96 : GEN_1028;
  assign GEN_1030 = 9'h61 == T_24222 ? T_18228_97 : GEN_1029;
  assign GEN_1031 = 9'h62 == T_24222 ? T_18228_98 : GEN_1030;
  assign GEN_1032 = 9'h63 == T_24222 ? T_18228_99 : GEN_1031;
  assign GEN_1033 = 9'h64 == T_24222 ? T_18228_100 : GEN_1032;
  assign GEN_1034 = 9'h65 == T_24222 ? T_18228_101 : GEN_1033;
  assign GEN_1035 = 9'h66 == T_24222 ? T_18228_102 : GEN_1034;
  assign GEN_1036 = 9'h67 == T_24222 ? T_18228_103 : GEN_1035;
  assign GEN_1037 = 9'h68 == T_24222 ? T_18228_104 : GEN_1036;
  assign GEN_1038 = 9'h69 == T_24222 ? T_18228_105 : GEN_1037;
  assign GEN_1039 = 9'h6a == T_24222 ? T_18228_106 : GEN_1038;
  assign GEN_1040 = 9'h6b == T_24222 ? T_18228_107 : GEN_1039;
  assign GEN_1041 = 9'h6c == T_24222 ? T_18228_108 : GEN_1040;
  assign GEN_1042 = 9'h6d == T_24222 ? T_18228_109 : GEN_1041;
  assign GEN_1043 = 9'h6e == T_24222 ? T_18228_110 : GEN_1042;
  assign GEN_1044 = 9'h6f == T_24222 ? T_18228_111 : GEN_1043;
  assign GEN_1045 = 9'h70 == T_24222 ? T_18228_112 : GEN_1044;
  assign GEN_1046 = 9'h71 == T_24222 ? T_18228_113 : GEN_1045;
  assign GEN_1047 = 9'h72 == T_24222 ? T_18228_114 : GEN_1046;
  assign GEN_1048 = 9'h73 == T_24222 ? T_18228_115 : GEN_1047;
  assign GEN_1049 = 9'h74 == T_24222 ? T_18228_116 : GEN_1048;
  assign GEN_1050 = 9'h75 == T_24222 ? T_18228_117 : GEN_1049;
  assign GEN_1051 = 9'h76 == T_24222 ? T_18228_118 : GEN_1050;
  assign GEN_1052 = 9'h77 == T_24222 ? T_18228_119 : GEN_1051;
  assign GEN_1053 = 9'h78 == T_24222 ? T_18228_120 : GEN_1052;
  assign GEN_1054 = 9'h79 == T_24222 ? T_18228_121 : GEN_1053;
  assign GEN_1055 = 9'h7a == T_24222 ? T_18228_122 : GEN_1054;
  assign GEN_1056 = 9'h7b == T_24222 ? T_18228_123 : GEN_1055;
  assign GEN_1057 = 9'h7c == T_24222 ? T_18228_124 : GEN_1056;
  assign GEN_1058 = 9'h7d == T_24222 ? T_18228_125 : GEN_1057;
  assign GEN_1059 = 9'h7e == T_24222 ? T_18228_126 : GEN_1058;
  assign GEN_1060 = 9'h7f == T_24222 ? T_18228_127 : GEN_1059;
  assign GEN_1061 = 9'h80 == T_24222 ? T_18228_128 : GEN_1060;
  assign GEN_1062 = 9'h81 == T_24222 ? T_18228_129 : GEN_1061;
  assign GEN_1063 = 9'h82 == T_24222 ? T_18228_130 : GEN_1062;
  assign GEN_1064 = 9'h83 == T_24222 ? T_18228_131 : GEN_1063;
  assign GEN_1065 = 9'h84 == T_24222 ? T_18228_132 : GEN_1064;
  assign GEN_1066 = 9'h85 == T_24222 ? T_18228_133 : GEN_1065;
  assign GEN_1067 = 9'h86 == T_24222 ? T_18228_134 : GEN_1066;
  assign GEN_1068 = 9'h87 == T_24222 ? T_18228_135 : GEN_1067;
  assign GEN_1069 = 9'h88 == T_24222 ? T_18228_136 : GEN_1068;
  assign GEN_1070 = 9'h89 == T_24222 ? T_18228_137 : GEN_1069;
  assign GEN_1071 = 9'h8a == T_24222 ? T_18228_138 : GEN_1070;
  assign GEN_1072 = 9'h8b == T_24222 ? T_18228_139 : GEN_1071;
  assign GEN_1073 = 9'h8c == T_24222 ? T_18228_140 : GEN_1072;
  assign GEN_1074 = 9'h8d == T_24222 ? T_18228_141 : GEN_1073;
  assign GEN_1075 = 9'h8e == T_24222 ? T_18228_142 : GEN_1074;
  assign GEN_1076 = 9'h8f == T_24222 ? T_18228_143 : GEN_1075;
  assign GEN_1077 = 9'h90 == T_24222 ? T_18228_144 : GEN_1076;
  assign GEN_1078 = 9'h91 == T_24222 ? T_18228_145 : GEN_1077;
  assign GEN_1079 = 9'h92 == T_24222 ? T_18228_146 : GEN_1078;
  assign GEN_1080 = 9'h93 == T_24222 ? T_18228_147 : GEN_1079;
  assign GEN_1081 = 9'h94 == T_24222 ? T_18228_148 : GEN_1080;
  assign GEN_1082 = 9'h95 == T_24222 ? T_18228_149 : GEN_1081;
  assign GEN_1083 = 9'h96 == T_24222 ? T_18228_150 : GEN_1082;
  assign GEN_1084 = 9'h97 == T_24222 ? T_18228_151 : GEN_1083;
  assign GEN_1085 = 9'h98 == T_24222 ? T_18228_152 : GEN_1084;
  assign GEN_1086 = 9'h99 == T_24222 ? T_18228_153 : GEN_1085;
  assign GEN_1087 = 9'h9a == T_24222 ? T_18228_154 : GEN_1086;
  assign GEN_1088 = 9'h9b == T_24222 ? T_18228_155 : GEN_1087;
  assign GEN_1089 = 9'h9c == T_24222 ? T_18228_156 : GEN_1088;
  assign GEN_1090 = 9'h9d == T_24222 ? T_18228_157 : GEN_1089;
  assign GEN_1091 = 9'h9e == T_24222 ? T_18228_158 : GEN_1090;
  assign GEN_1092 = 9'h9f == T_24222 ? T_18228_159 : GEN_1091;
  assign GEN_1093 = 9'ha0 == T_24222 ? T_18228_160 : GEN_1092;
  assign GEN_1094 = 9'ha1 == T_24222 ? T_18228_161 : GEN_1093;
  assign GEN_1095 = 9'ha2 == T_24222 ? T_18228_162 : GEN_1094;
  assign GEN_1096 = 9'ha3 == T_24222 ? T_18228_163 : GEN_1095;
  assign GEN_1097 = 9'ha4 == T_24222 ? T_18228_164 : GEN_1096;
  assign GEN_1098 = 9'ha5 == T_24222 ? T_18228_165 : GEN_1097;
  assign GEN_1099 = 9'ha6 == T_24222 ? T_18228_166 : GEN_1098;
  assign GEN_1100 = 9'ha7 == T_24222 ? T_18228_167 : GEN_1099;
  assign GEN_1101 = 9'ha8 == T_24222 ? T_18228_168 : GEN_1100;
  assign GEN_1102 = 9'ha9 == T_24222 ? T_18228_169 : GEN_1101;
  assign GEN_1103 = 9'haa == T_24222 ? T_18228_170 : GEN_1102;
  assign GEN_1104 = 9'hab == T_24222 ? T_18228_171 : GEN_1103;
  assign GEN_1105 = 9'hac == T_24222 ? T_18228_172 : GEN_1104;
  assign GEN_1106 = 9'had == T_24222 ? T_18228_173 : GEN_1105;
  assign GEN_1107 = 9'hae == T_24222 ? T_18228_174 : GEN_1106;
  assign GEN_1108 = 9'haf == T_24222 ? T_18228_175 : GEN_1107;
  assign GEN_1109 = 9'hb0 == T_24222 ? T_18228_176 : GEN_1108;
  assign GEN_1110 = 9'hb1 == T_24222 ? T_18228_177 : GEN_1109;
  assign GEN_1111 = 9'hb2 == T_24222 ? T_18228_178 : GEN_1110;
  assign GEN_1112 = 9'hb3 == T_24222 ? T_18228_179 : GEN_1111;
  assign GEN_1113 = 9'hb4 == T_24222 ? T_18228_180 : GEN_1112;
  assign GEN_1114 = 9'hb5 == T_24222 ? T_18228_181 : GEN_1113;
  assign GEN_1115 = 9'hb6 == T_24222 ? T_18228_182 : GEN_1114;
  assign GEN_1116 = 9'hb7 == T_24222 ? T_18228_183 : GEN_1115;
  assign GEN_1117 = 9'hb8 == T_24222 ? T_18228_184 : GEN_1116;
  assign GEN_1118 = 9'hb9 == T_24222 ? T_18228_185 : GEN_1117;
  assign GEN_1119 = 9'hba == T_24222 ? T_18228_186 : GEN_1118;
  assign GEN_1120 = 9'hbb == T_24222 ? T_18228_187 : GEN_1119;
  assign GEN_1121 = 9'hbc == T_24222 ? T_18228_188 : GEN_1120;
  assign GEN_1122 = 9'hbd == T_24222 ? T_18228_189 : GEN_1121;
  assign GEN_1123 = 9'hbe == T_24222 ? T_18228_190 : GEN_1122;
  assign GEN_1124 = 9'hbf == T_24222 ? T_18228_191 : GEN_1123;
  assign GEN_1125 = 9'hc0 == T_24222 ? T_18228_192 : GEN_1124;
  assign GEN_1126 = 9'hc1 == T_24222 ? T_18228_193 : GEN_1125;
  assign GEN_1127 = 9'hc2 == T_24222 ? T_18228_194 : GEN_1126;
  assign GEN_1128 = 9'hc3 == T_24222 ? T_18228_195 : GEN_1127;
  assign GEN_1129 = 9'hc4 == T_24222 ? T_18228_196 : GEN_1128;
  assign GEN_1130 = 9'hc5 == T_24222 ? T_18228_197 : GEN_1129;
  assign GEN_1131 = 9'hc6 == T_24222 ? T_18228_198 : GEN_1130;
  assign GEN_1132 = 9'hc7 == T_24222 ? T_18228_199 : GEN_1131;
  assign GEN_1133 = 9'hc8 == T_24222 ? T_18228_200 : GEN_1132;
  assign GEN_1134 = 9'hc9 == T_24222 ? T_18228_201 : GEN_1133;
  assign GEN_1135 = 9'hca == T_24222 ? T_18228_202 : GEN_1134;
  assign GEN_1136 = 9'hcb == T_24222 ? T_18228_203 : GEN_1135;
  assign GEN_1137 = 9'hcc == T_24222 ? T_18228_204 : GEN_1136;
  assign GEN_1138 = 9'hcd == T_24222 ? T_18228_205 : GEN_1137;
  assign GEN_1139 = 9'hce == T_24222 ? T_18228_206 : GEN_1138;
  assign GEN_1140 = 9'hcf == T_24222 ? T_18228_207 : GEN_1139;
  assign GEN_1141 = 9'hd0 == T_24222 ? T_18228_208 : GEN_1140;
  assign GEN_1142 = 9'hd1 == T_24222 ? T_18228_209 : GEN_1141;
  assign GEN_1143 = 9'hd2 == T_24222 ? T_18228_210 : GEN_1142;
  assign GEN_1144 = 9'hd3 == T_24222 ? T_18228_211 : GEN_1143;
  assign GEN_1145 = 9'hd4 == T_24222 ? T_18228_212 : GEN_1144;
  assign GEN_1146 = 9'hd5 == T_24222 ? T_18228_213 : GEN_1145;
  assign GEN_1147 = 9'hd6 == T_24222 ? T_18228_214 : GEN_1146;
  assign GEN_1148 = 9'hd7 == T_24222 ? T_18228_215 : GEN_1147;
  assign GEN_1149 = 9'hd8 == T_24222 ? T_18228_216 : GEN_1148;
  assign GEN_1150 = 9'hd9 == T_24222 ? T_18228_217 : GEN_1149;
  assign GEN_1151 = 9'hda == T_24222 ? T_18228_218 : GEN_1150;
  assign GEN_1152 = 9'hdb == T_24222 ? T_18228_219 : GEN_1151;
  assign GEN_1153 = 9'hdc == T_24222 ? T_18228_220 : GEN_1152;
  assign GEN_1154 = 9'hdd == T_24222 ? T_18228_221 : GEN_1153;
  assign GEN_1155 = 9'hde == T_24222 ? T_18228_222 : GEN_1154;
  assign GEN_1156 = 9'hdf == T_24222 ? T_18228_223 : GEN_1155;
  assign GEN_1157 = 9'he0 == T_24222 ? T_18228_224 : GEN_1156;
  assign GEN_1158 = 9'he1 == T_24222 ? T_18228_225 : GEN_1157;
  assign GEN_1159 = 9'he2 == T_24222 ? T_18228_226 : GEN_1158;
  assign GEN_1160 = 9'he3 == T_24222 ? T_18228_227 : GEN_1159;
  assign GEN_1161 = 9'he4 == T_24222 ? T_18228_228 : GEN_1160;
  assign GEN_1162 = 9'he5 == T_24222 ? T_18228_229 : GEN_1161;
  assign GEN_1163 = 9'he6 == T_24222 ? T_18228_230 : GEN_1162;
  assign GEN_1164 = 9'he7 == T_24222 ? T_18228_231 : GEN_1163;
  assign GEN_1165 = 9'he8 == T_24222 ? T_18228_232 : GEN_1164;
  assign GEN_1166 = 9'he9 == T_24222 ? T_18228_233 : GEN_1165;
  assign GEN_1167 = 9'hea == T_24222 ? T_18228_234 : GEN_1166;
  assign GEN_1168 = 9'heb == T_24222 ? T_18228_235 : GEN_1167;
  assign GEN_1169 = 9'hec == T_24222 ? T_18228_236 : GEN_1168;
  assign GEN_1170 = 9'hed == T_24222 ? T_18228_237 : GEN_1169;
  assign GEN_1171 = 9'hee == T_24222 ? T_18228_238 : GEN_1170;
  assign GEN_1172 = 9'hef == T_24222 ? T_18228_239 : GEN_1171;
  assign GEN_1173 = 9'hf0 == T_24222 ? T_18228_240 : GEN_1172;
  assign GEN_1174 = 9'hf1 == T_24222 ? T_18228_241 : GEN_1173;
  assign GEN_1175 = 9'hf2 == T_24222 ? T_18228_242 : GEN_1174;
  assign GEN_1176 = 9'hf3 == T_24222 ? T_18228_243 : GEN_1175;
  assign GEN_1177 = 9'hf4 == T_24222 ? T_18228_244 : GEN_1176;
  assign GEN_1178 = 9'hf5 == T_24222 ? T_18228_245 : GEN_1177;
  assign GEN_1179 = 9'hf6 == T_24222 ? T_18228_246 : GEN_1178;
  assign GEN_1180 = 9'hf7 == T_24222 ? T_18228_247 : GEN_1179;
  assign GEN_1181 = 9'hf8 == T_24222 ? T_18228_248 : GEN_1180;
  assign GEN_1182 = 9'hf9 == T_24222 ? T_18228_249 : GEN_1181;
  assign GEN_1183 = 9'hfa == T_24222 ? T_18228_250 : GEN_1182;
  assign GEN_1184 = 9'hfb == T_24222 ? T_18228_251 : GEN_1183;
  assign GEN_1185 = 9'hfc == T_24222 ? T_18228_252 : GEN_1184;
  assign GEN_1186 = 9'hfd == T_24222 ? T_18228_253 : GEN_1185;
  assign GEN_1187 = 9'hfe == T_24222 ? T_18228_254 : GEN_1186;
  assign GEN_1188 = 9'hff == T_24222 ? T_18228_255 : GEN_1187;
  assign GEN_1189 = 9'h100 == T_24222 ? T_18228_256 : GEN_1188;
  assign GEN_1190 = 9'h101 == T_24222 ? T_18228_257 : GEN_1189;
  assign GEN_1191 = 9'h102 == T_24222 ? T_18228_258 : GEN_1190;
  assign GEN_1192 = 9'h103 == T_24222 ? T_18228_259 : GEN_1191;
  assign GEN_1193 = 9'h104 == T_24222 ? T_18228_260 : GEN_1192;
  assign GEN_1194 = 9'h105 == T_24222 ? T_18228_261 : GEN_1193;
  assign GEN_1195 = 9'h106 == T_24222 ? T_18228_262 : GEN_1194;
  assign GEN_1196 = 9'h107 == T_24222 ? T_18228_263 : GEN_1195;
  assign GEN_1197 = 9'h108 == T_24222 ? T_18228_264 : GEN_1196;
  assign GEN_1198 = 9'h109 == T_24222 ? T_18228_265 : GEN_1197;
  assign GEN_1199 = 9'h10a == T_24222 ? T_18228_266 : GEN_1198;
  assign GEN_1200 = 9'h10b == T_24222 ? T_18228_267 : GEN_1199;
  assign GEN_1201 = 9'h10c == T_24222 ? T_18228_268 : GEN_1200;
  assign GEN_1202 = 9'h10d == T_24222 ? T_18228_269 : GEN_1201;
  assign GEN_1203 = 9'h10e == T_24222 ? T_18228_270 : GEN_1202;
  assign GEN_1204 = 9'h10f == T_24222 ? T_18228_271 : GEN_1203;
  assign GEN_1205 = 9'h110 == T_24222 ? T_18228_272 : GEN_1204;
  assign GEN_1206 = 9'h111 == T_24222 ? T_18228_273 : GEN_1205;
  assign GEN_1207 = 9'h112 == T_24222 ? T_18228_274 : GEN_1206;
  assign GEN_1208 = 9'h113 == T_24222 ? T_18228_275 : GEN_1207;
  assign GEN_1209 = 9'h114 == T_24222 ? T_18228_276 : GEN_1208;
  assign GEN_1210 = 9'h115 == T_24222 ? T_18228_277 : GEN_1209;
  assign GEN_1211 = 9'h116 == T_24222 ? T_18228_278 : GEN_1210;
  assign GEN_1212 = 9'h117 == T_24222 ? T_18228_279 : GEN_1211;
  assign GEN_1213 = 9'h118 == T_24222 ? T_18228_280 : GEN_1212;
  assign GEN_1214 = 9'h119 == T_24222 ? T_18228_281 : GEN_1213;
  assign GEN_1215 = 9'h11a == T_24222 ? T_18228_282 : GEN_1214;
  assign GEN_1216 = 9'h11b == T_24222 ? T_18228_283 : GEN_1215;
  assign GEN_1217 = 9'h11c == T_24222 ? T_18228_284 : GEN_1216;
  assign GEN_1218 = 9'h11d == T_24222 ? T_18228_285 : GEN_1217;
  assign GEN_1219 = 9'h11e == T_24222 ? T_18228_286 : GEN_1218;
  assign GEN_1220 = 9'h11f == T_24222 ? T_18228_287 : GEN_1219;
  assign GEN_1221 = 9'h120 == T_24222 ? T_18228_288 : GEN_1220;
  assign GEN_1222 = 9'h121 == T_24222 ? T_18228_289 : GEN_1221;
  assign GEN_1223 = 9'h122 == T_24222 ? T_18228_290 : GEN_1222;
  assign GEN_1224 = 9'h123 == T_24222 ? T_18228_291 : GEN_1223;
  assign GEN_1225 = 9'h124 == T_24222 ? T_18228_292 : GEN_1224;
  assign GEN_1226 = 9'h125 == T_24222 ? T_18228_293 : GEN_1225;
  assign GEN_1227 = 9'h126 == T_24222 ? T_18228_294 : GEN_1226;
  assign GEN_1228 = 9'h127 == T_24222 ? T_18228_295 : GEN_1227;
  assign GEN_1229 = 9'h128 == T_24222 ? T_18228_296 : GEN_1228;
  assign GEN_1230 = 9'h129 == T_24222 ? T_18228_297 : GEN_1229;
  assign GEN_1231 = 9'h12a == T_24222 ? T_18228_298 : GEN_1230;
  assign GEN_1232 = 9'h12b == T_24222 ? T_18228_299 : GEN_1231;
  assign GEN_1233 = 9'h12c == T_24222 ? T_18228_300 : GEN_1232;
  assign GEN_1234 = 9'h12d == T_24222 ? T_18228_301 : GEN_1233;
  assign GEN_1235 = 9'h12e == T_24222 ? T_18228_302 : GEN_1234;
  assign GEN_1236 = 9'h12f == T_24222 ? T_18228_303 : GEN_1235;
  assign GEN_1237 = 9'h130 == T_24222 ? T_18228_304 : GEN_1236;
  assign GEN_1238 = 9'h131 == T_24222 ? T_18228_305 : GEN_1237;
  assign GEN_1239 = 9'h132 == T_24222 ? T_18228_306 : GEN_1238;
  assign GEN_1240 = 9'h133 == T_24222 ? T_18228_307 : GEN_1239;
  assign GEN_1241 = 9'h134 == T_24222 ? T_18228_308 : GEN_1240;
  assign GEN_1242 = 9'h135 == T_24222 ? T_18228_309 : GEN_1241;
  assign GEN_1243 = 9'h136 == T_24222 ? T_18228_310 : GEN_1242;
  assign GEN_1244 = 9'h137 == T_24222 ? T_18228_311 : GEN_1243;
  assign GEN_1245 = 9'h138 == T_24222 ? T_18228_312 : GEN_1244;
  assign GEN_1246 = 9'h139 == T_24222 ? T_18228_313 : GEN_1245;
  assign GEN_1247 = 9'h13a == T_24222 ? T_18228_314 : GEN_1246;
  assign GEN_1248 = 9'h13b == T_24222 ? T_18228_315 : GEN_1247;
  assign GEN_1249 = 9'h13c == T_24222 ? T_18228_316 : GEN_1248;
  assign GEN_1250 = 9'h13d == T_24222 ? T_18228_317 : GEN_1249;
  assign GEN_1251 = 9'h13e == T_24222 ? T_18228_318 : GEN_1250;
  assign GEN_1252 = 9'h13f == T_24222 ? T_18228_319 : GEN_1251;
  assign GEN_1253 = 9'h140 == T_24222 ? T_18228_320 : GEN_1252;
  assign GEN_1254 = 9'h141 == T_24222 ? T_18228_321 : GEN_1253;
  assign GEN_1255 = 9'h142 == T_24222 ? T_18228_322 : GEN_1254;
  assign GEN_1256 = 9'h143 == T_24222 ? T_18228_323 : GEN_1255;
  assign GEN_1257 = 9'h144 == T_24222 ? T_18228_324 : GEN_1256;
  assign GEN_1258 = 9'h145 == T_24222 ? T_18228_325 : GEN_1257;
  assign GEN_1259 = 9'h146 == T_24222 ? T_18228_326 : GEN_1258;
  assign GEN_1260 = 9'h147 == T_24222 ? T_18228_327 : GEN_1259;
  assign GEN_1261 = 9'h148 == T_24222 ? T_18228_328 : GEN_1260;
  assign GEN_1262 = 9'h149 == T_24222 ? T_18228_329 : GEN_1261;
  assign GEN_1263 = 9'h14a == T_24222 ? T_18228_330 : GEN_1262;
  assign GEN_1264 = 9'h14b == T_24222 ? T_18228_331 : GEN_1263;
  assign GEN_1265 = 9'h14c == T_24222 ? T_18228_332 : GEN_1264;
  assign GEN_1266 = 9'h14d == T_24222 ? T_18228_333 : GEN_1265;
  assign GEN_1267 = 9'h14e == T_24222 ? T_18228_334 : GEN_1266;
  assign GEN_1268 = 9'h14f == T_24222 ? T_18228_335 : GEN_1267;
  assign GEN_1269 = 9'h150 == T_24222 ? T_18228_336 : GEN_1268;
  assign GEN_1270 = 9'h151 == T_24222 ? T_18228_337 : GEN_1269;
  assign GEN_1271 = 9'h152 == T_24222 ? T_18228_338 : GEN_1270;
  assign GEN_1272 = 9'h153 == T_24222 ? T_18228_339 : GEN_1271;
  assign GEN_1273 = 9'h154 == T_24222 ? T_18228_340 : GEN_1272;
  assign GEN_1274 = 9'h155 == T_24222 ? T_18228_341 : GEN_1273;
  assign GEN_1275 = 9'h156 == T_24222 ? T_18228_342 : GEN_1274;
  assign GEN_1276 = 9'h157 == T_24222 ? T_18228_343 : GEN_1275;
  assign GEN_1277 = 9'h158 == T_24222 ? T_18228_344 : GEN_1276;
  assign GEN_1278 = 9'h159 == T_24222 ? T_18228_345 : GEN_1277;
  assign GEN_1279 = 9'h15a == T_24222 ? T_18228_346 : GEN_1278;
  assign GEN_1280 = 9'h15b == T_24222 ? T_18228_347 : GEN_1279;
  assign GEN_1281 = 9'h15c == T_24222 ? T_18228_348 : GEN_1280;
  assign GEN_1282 = 9'h15d == T_24222 ? T_18228_349 : GEN_1281;
  assign GEN_1283 = 9'h15e == T_24222 ? T_18228_350 : GEN_1282;
  assign GEN_1284 = 9'h15f == T_24222 ? T_18228_351 : GEN_1283;
  assign GEN_1285 = 9'h160 == T_24222 ? T_18228_352 : GEN_1284;
  assign GEN_1286 = 9'h161 == T_24222 ? T_18228_353 : GEN_1285;
  assign GEN_1287 = 9'h162 == T_24222 ? T_18228_354 : GEN_1286;
  assign GEN_1288 = 9'h163 == T_24222 ? T_18228_355 : GEN_1287;
  assign GEN_1289 = 9'h164 == T_24222 ? T_18228_356 : GEN_1288;
  assign GEN_1290 = 9'h165 == T_24222 ? T_18228_357 : GEN_1289;
  assign GEN_1291 = 9'h166 == T_24222 ? T_18228_358 : GEN_1290;
  assign GEN_1292 = 9'h167 == T_24222 ? T_18228_359 : GEN_1291;
  assign GEN_1293 = 9'h168 == T_24222 ? T_18228_360 : GEN_1292;
  assign GEN_1294 = 9'h169 == T_24222 ? T_18228_361 : GEN_1293;
  assign GEN_1295 = 9'h16a == T_24222 ? T_18228_362 : GEN_1294;
  assign GEN_1296 = 9'h16b == T_24222 ? T_18228_363 : GEN_1295;
  assign GEN_1297 = 9'h16c == T_24222 ? T_18228_364 : GEN_1296;
  assign GEN_1298 = 9'h16d == T_24222 ? T_18228_365 : GEN_1297;
  assign GEN_1299 = 9'h16e == T_24222 ? T_18228_366 : GEN_1298;
  assign GEN_1300 = 9'h16f == T_24222 ? T_18228_367 : GEN_1299;
  assign GEN_1301 = 9'h170 == T_24222 ? T_18228_368 : GEN_1300;
  assign GEN_1302 = 9'h171 == T_24222 ? T_18228_369 : GEN_1301;
  assign GEN_1303 = 9'h172 == T_24222 ? T_18228_370 : GEN_1302;
  assign GEN_1304 = 9'h173 == T_24222 ? T_18228_371 : GEN_1303;
  assign GEN_1305 = 9'h174 == T_24222 ? T_18228_372 : GEN_1304;
  assign GEN_1306 = 9'h175 == T_24222 ? T_18228_373 : GEN_1305;
  assign GEN_1307 = 9'h176 == T_24222 ? T_18228_374 : GEN_1306;
  assign GEN_1308 = 9'h177 == T_24222 ? T_18228_375 : GEN_1307;
  assign GEN_1309 = 9'h178 == T_24222 ? T_18228_376 : GEN_1308;
  assign GEN_1310 = 9'h179 == T_24222 ? T_18228_377 : GEN_1309;
  assign GEN_1311 = 9'h17a == T_24222 ? T_18228_378 : GEN_1310;
  assign GEN_1312 = 9'h17b == T_24222 ? T_18228_379 : GEN_1311;
  assign GEN_1313 = 9'h17c == T_24222 ? T_18228_380 : GEN_1312;
  assign GEN_1314 = 9'h17d == T_24222 ? T_18228_381 : GEN_1313;
  assign GEN_1315 = 9'h17e == T_24222 ? T_18228_382 : GEN_1314;
  assign GEN_1316 = 9'h17f == T_24222 ? T_18228_383 : GEN_1315;
  assign GEN_1317 = 9'h180 == T_24222 ? T_18228_384 : GEN_1316;
  assign GEN_1318 = 9'h181 == T_24222 ? T_18228_385 : GEN_1317;
  assign GEN_1319 = 9'h182 == T_24222 ? T_18228_386 : GEN_1318;
  assign GEN_1320 = 9'h183 == T_24222 ? T_18228_387 : GEN_1319;
  assign GEN_1321 = 9'h184 == T_24222 ? T_18228_388 : GEN_1320;
  assign GEN_1322 = 9'h185 == T_24222 ? T_18228_389 : GEN_1321;
  assign GEN_1323 = 9'h186 == T_24222 ? T_18228_390 : GEN_1322;
  assign GEN_1324 = 9'h187 == T_24222 ? T_18228_391 : GEN_1323;
  assign GEN_1325 = 9'h188 == T_24222 ? T_18228_392 : GEN_1324;
  assign GEN_1326 = 9'h189 == T_24222 ? T_18228_393 : GEN_1325;
  assign GEN_1327 = 9'h18a == T_24222 ? T_18228_394 : GEN_1326;
  assign GEN_1328 = 9'h18b == T_24222 ? T_18228_395 : GEN_1327;
  assign GEN_1329 = 9'h18c == T_24222 ? T_18228_396 : GEN_1328;
  assign GEN_1330 = 9'h18d == T_24222 ? T_18228_397 : GEN_1329;
  assign GEN_1331 = 9'h18e == T_24222 ? T_18228_398 : GEN_1330;
  assign GEN_1332 = 9'h18f == T_24222 ? T_18228_399 : GEN_1331;
  assign GEN_1333 = 9'h190 == T_24222 ? T_18228_400 : GEN_1332;
  assign GEN_1334 = 9'h191 == T_24222 ? T_18228_401 : GEN_1333;
  assign GEN_1335 = 9'h192 == T_24222 ? T_18228_402 : GEN_1334;
  assign GEN_1336 = 9'h193 == T_24222 ? T_18228_403 : GEN_1335;
  assign GEN_1337 = 9'h194 == T_24222 ? T_18228_404 : GEN_1336;
  assign GEN_1338 = 9'h195 == T_24222 ? T_18228_405 : GEN_1337;
  assign GEN_1339 = 9'h196 == T_24222 ? T_18228_406 : GEN_1338;
  assign GEN_1340 = 9'h197 == T_24222 ? T_18228_407 : GEN_1339;
  assign GEN_1341 = 9'h198 == T_24222 ? T_18228_408 : GEN_1340;
  assign GEN_1342 = 9'h199 == T_24222 ? T_18228_409 : GEN_1341;
  assign GEN_1343 = 9'h19a == T_24222 ? T_18228_410 : GEN_1342;
  assign GEN_1344 = 9'h19b == T_24222 ? T_18228_411 : GEN_1343;
  assign GEN_1345 = 9'h19c == T_24222 ? T_18228_412 : GEN_1344;
  assign GEN_1346 = 9'h19d == T_24222 ? T_18228_413 : GEN_1345;
  assign GEN_1347 = 9'h19e == T_24222 ? T_18228_414 : GEN_1346;
  assign GEN_1348 = 9'h19f == T_24222 ? T_18228_415 : GEN_1347;
  assign GEN_1349 = 9'h1a0 == T_24222 ? T_18228_416 : GEN_1348;
  assign GEN_1350 = 9'h1a1 == T_24222 ? T_18228_417 : GEN_1349;
  assign GEN_1351 = 9'h1a2 == T_24222 ? T_18228_418 : GEN_1350;
  assign GEN_1352 = 9'h1a3 == T_24222 ? T_18228_419 : GEN_1351;
  assign GEN_1353 = 9'h1a4 == T_24222 ? T_18228_420 : GEN_1352;
  assign GEN_1354 = 9'h1a5 == T_24222 ? T_18228_421 : GEN_1353;
  assign GEN_1355 = 9'h1a6 == T_24222 ? T_18228_422 : GEN_1354;
  assign GEN_1356 = 9'h1a7 == T_24222 ? T_18228_423 : GEN_1355;
  assign GEN_1357 = 9'h1a8 == T_24222 ? T_18228_424 : GEN_1356;
  assign GEN_1358 = 9'h1a9 == T_24222 ? T_18228_425 : GEN_1357;
  assign GEN_1359 = 9'h1aa == T_24222 ? T_18228_426 : GEN_1358;
  assign GEN_1360 = 9'h1ab == T_24222 ? T_18228_427 : GEN_1359;
  assign GEN_1361 = 9'h1ac == T_24222 ? T_18228_428 : GEN_1360;
  assign GEN_1362 = 9'h1ad == T_24222 ? T_18228_429 : GEN_1361;
  assign GEN_1363 = 9'h1ae == T_24222 ? T_18228_430 : GEN_1362;
  assign GEN_1364 = 9'h1af == T_24222 ? T_18228_431 : GEN_1363;
  assign GEN_1365 = 9'h1b0 == T_24222 ? T_18228_432 : GEN_1364;
  assign GEN_1366 = 9'h1b1 == T_24222 ? T_18228_433 : GEN_1365;
  assign GEN_1367 = 9'h1b2 == T_24222 ? T_18228_434 : GEN_1366;
  assign GEN_1368 = 9'h1b3 == T_24222 ? T_18228_435 : GEN_1367;
  assign GEN_1369 = 9'h1b4 == T_24222 ? T_18228_436 : GEN_1368;
  assign GEN_1370 = 9'h1b5 == T_24222 ? T_18228_437 : GEN_1369;
  assign GEN_1371 = 9'h1b6 == T_24222 ? T_18228_438 : GEN_1370;
  assign GEN_1372 = 9'h1b7 == T_24222 ? T_18228_439 : GEN_1371;
  assign GEN_1373 = 9'h1b8 == T_24222 ? T_18228_440 : GEN_1372;
  assign GEN_1374 = 9'h1b9 == T_24222 ? T_18228_441 : GEN_1373;
  assign GEN_1375 = 9'h1ba == T_24222 ? T_18228_442 : GEN_1374;
  assign GEN_1376 = 9'h1bb == T_24222 ? T_18228_443 : GEN_1375;
  assign GEN_1377 = 9'h1bc == T_24222 ? T_18228_444 : GEN_1376;
  assign GEN_1378 = 9'h1bd == T_24222 ? T_18228_445 : GEN_1377;
  assign GEN_1379 = 9'h1be == T_24222 ? T_18228_446 : GEN_1378;
  assign GEN_1380 = 9'h1bf == T_24222 ? T_18228_447 : GEN_1379;
  assign GEN_1381 = 9'h1c0 == T_24222 ? T_18228_448 : GEN_1380;
  assign GEN_1382 = 9'h1c1 == T_24222 ? T_18228_449 : GEN_1381;
  assign GEN_1383 = 9'h1c2 == T_24222 ? T_18228_450 : GEN_1382;
  assign GEN_1384 = 9'h1c3 == T_24222 ? T_18228_451 : GEN_1383;
  assign GEN_1385 = 9'h1c4 == T_24222 ? T_18228_452 : GEN_1384;
  assign GEN_1386 = 9'h1c5 == T_24222 ? T_18228_453 : GEN_1385;
  assign GEN_1387 = 9'h1c6 == T_24222 ? T_18228_454 : GEN_1386;
  assign GEN_1388 = 9'h1c7 == T_24222 ? T_18228_455 : GEN_1387;
  assign GEN_1389 = 9'h1c8 == T_24222 ? T_18228_456 : GEN_1388;
  assign GEN_1390 = 9'h1c9 == T_24222 ? T_18228_457 : GEN_1389;
  assign GEN_1391 = 9'h1ca == T_24222 ? T_18228_458 : GEN_1390;
  assign GEN_1392 = 9'h1cb == T_24222 ? T_18228_459 : GEN_1391;
  assign GEN_1393 = 9'h1cc == T_24222 ? T_18228_460 : GEN_1392;
  assign GEN_1394 = 9'h1cd == T_24222 ? T_18228_461 : GEN_1393;
  assign GEN_1395 = 9'h1ce == T_24222 ? T_18228_462 : GEN_1394;
  assign GEN_1396 = 9'h1cf == T_24222 ? T_18228_463 : GEN_1395;
  assign GEN_1397 = 9'h1d0 == T_24222 ? T_18228_464 : GEN_1396;
  assign GEN_1398 = 9'h1d1 == T_24222 ? T_18228_465 : GEN_1397;
  assign GEN_1399 = 9'h1d2 == T_24222 ? T_18228_466 : GEN_1398;
  assign GEN_1400 = 9'h1d3 == T_24222 ? T_18228_467 : GEN_1399;
  assign GEN_1401 = 9'h1d4 == T_24222 ? T_18228_468 : GEN_1400;
  assign GEN_1402 = 9'h1d5 == T_24222 ? T_18228_469 : GEN_1401;
  assign GEN_1403 = 9'h1d6 == T_24222 ? T_18228_470 : GEN_1402;
  assign GEN_1404 = 9'h1d7 == T_24222 ? T_18228_471 : GEN_1403;
  assign GEN_1405 = 9'h1d8 == T_24222 ? T_18228_472 : GEN_1404;
  assign GEN_1406 = 9'h1d9 == T_24222 ? T_18228_473 : GEN_1405;
  assign GEN_1407 = 9'h1da == T_24222 ? T_18228_474 : GEN_1406;
  assign GEN_1408 = 9'h1db == T_24222 ? T_18228_475 : GEN_1407;
  assign GEN_1409 = 9'h1dc == T_24222 ? T_18228_476 : GEN_1408;
  assign GEN_1410 = 9'h1dd == T_24222 ? T_18228_477 : GEN_1409;
  assign GEN_1411 = 9'h1de == T_24222 ? T_18228_478 : GEN_1410;
  assign GEN_1412 = 9'h1df == T_24222 ? T_18228_479 : GEN_1411;
  assign GEN_1413 = 9'h1e0 == T_24222 ? T_18228_480 : GEN_1412;
  assign GEN_1414 = 9'h1e1 == T_24222 ? T_18228_481 : GEN_1413;
  assign GEN_1415 = 9'h1e2 == T_24222 ? T_18228_482 : GEN_1414;
  assign GEN_1416 = 9'h1e3 == T_24222 ? T_18228_483 : GEN_1415;
  assign GEN_1417 = 9'h1e4 == T_24222 ? T_18228_484 : GEN_1416;
  assign GEN_1418 = 9'h1e5 == T_24222 ? T_18228_485 : GEN_1417;
  assign GEN_1419 = 9'h1e6 == T_24222 ? T_18228_486 : GEN_1418;
  assign GEN_1420 = 9'h1e7 == T_24222 ? T_18228_487 : GEN_1419;
  assign GEN_1421 = 9'h1e8 == T_24222 ? T_18228_488 : GEN_1420;
  assign GEN_1422 = 9'h1e9 == T_24222 ? T_18228_489 : GEN_1421;
  assign GEN_1423 = 9'h1ea == T_24222 ? T_18228_490 : GEN_1422;
  assign GEN_1424 = 9'h1eb == T_24222 ? T_18228_491 : GEN_1423;
  assign GEN_1425 = 9'h1ec == T_24222 ? T_18228_492 : GEN_1424;
  assign GEN_1426 = 9'h1ed == T_24222 ? T_18228_493 : GEN_1425;
  assign GEN_1427 = 9'h1ee == T_24222 ? T_18228_494 : GEN_1426;
  assign GEN_1428 = 9'h1ef == T_24222 ? T_18228_495 : GEN_1427;
  assign GEN_1429 = 9'h1f0 == T_24222 ? T_18228_496 : GEN_1428;
  assign GEN_1430 = 9'h1f1 == T_24222 ? T_18228_497 : GEN_1429;
  assign GEN_1431 = 9'h1f2 == T_24222 ? T_18228_498 : GEN_1430;
  assign GEN_1432 = 9'h1f3 == T_24222 ? T_18228_499 : GEN_1431;
  assign GEN_1433 = 9'h1f4 == T_24222 ? T_18228_500 : GEN_1432;
  assign GEN_1434 = 9'h1f5 == T_24222 ? T_18228_501 : GEN_1433;
  assign GEN_1435 = 9'h1f6 == T_24222 ? T_18228_502 : GEN_1434;
  assign GEN_1436 = 9'h1f7 == T_24222 ? T_18228_503 : GEN_1435;
  assign GEN_1437 = 9'h1f8 == T_24222 ? T_18228_504 : GEN_1436;
  assign GEN_1438 = 9'h1f9 == T_24222 ? T_18228_505 : GEN_1437;
  assign GEN_1439 = 9'h1fa == T_24222 ? T_18228_506 : GEN_1438;
  assign GEN_1440 = 9'h1fb == T_24222 ? T_18228_507 : GEN_1439;
  assign GEN_1441 = 9'h1fc == T_24222 ? T_18228_508 : GEN_1440;
  assign GEN_1442 = 9'h1fd == T_24222 ? T_18228_509 : GEN_1441;
  assign GEN_1443 = 9'h1fe == T_24222 ? T_18228_510 : GEN_1442;
  assign GEN_1444 = 9'h1ff == T_24222 ? T_18228_511 : GEN_1443;
  assign T_24257 = T_3205_bits_read ? GEN_3 : GEN_4;
  assign GEN_5 = GEN_1955;
  assign GEN_1445 = 9'h1 == T_24222 ? T_20952_1 : T_20952_0;
  assign GEN_1446 = 9'h2 == T_24222 ? T_20952_2 : GEN_1445;
  assign GEN_1447 = 9'h3 == T_24222 ? T_20952_3 : GEN_1446;
  assign GEN_1448 = 9'h4 == T_24222 ? T_20952_4 : GEN_1447;
  assign GEN_1449 = 9'h5 == T_24222 ? T_20952_5 : GEN_1448;
  assign GEN_1450 = 9'h6 == T_24222 ? T_20952_6 : GEN_1449;
  assign GEN_1451 = 9'h7 == T_24222 ? T_20952_7 : GEN_1450;
  assign GEN_1452 = 9'h8 == T_24222 ? T_20952_8 : GEN_1451;
  assign GEN_1453 = 9'h9 == T_24222 ? T_20952_9 : GEN_1452;
  assign GEN_1454 = 9'ha == T_24222 ? T_20952_10 : GEN_1453;
  assign GEN_1455 = 9'hb == T_24222 ? T_20952_11 : GEN_1454;
  assign GEN_1456 = 9'hc == T_24222 ? T_20952_12 : GEN_1455;
  assign GEN_1457 = 9'hd == T_24222 ? T_20952_13 : GEN_1456;
  assign GEN_1458 = 9'he == T_24222 ? T_20952_14 : GEN_1457;
  assign GEN_1459 = 9'hf == T_24222 ? T_20952_15 : GEN_1458;
  assign GEN_1460 = 9'h10 == T_24222 ? T_20952_16 : GEN_1459;
  assign GEN_1461 = 9'h11 == T_24222 ? T_20952_17 : GEN_1460;
  assign GEN_1462 = 9'h12 == T_24222 ? T_20952_18 : GEN_1461;
  assign GEN_1463 = 9'h13 == T_24222 ? T_20952_19 : GEN_1462;
  assign GEN_1464 = 9'h14 == T_24222 ? T_20952_20 : GEN_1463;
  assign GEN_1465 = 9'h15 == T_24222 ? T_20952_21 : GEN_1464;
  assign GEN_1466 = 9'h16 == T_24222 ? T_20952_22 : GEN_1465;
  assign GEN_1467 = 9'h17 == T_24222 ? T_20952_23 : GEN_1466;
  assign GEN_1468 = 9'h18 == T_24222 ? T_20952_24 : GEN_1467;
  assign GEN_1469 = 9'h19 == T_24222 ? T_20952_25 : GEN_1468;
  assign GEN_1470 = 9'h1a == T_24222 ? T_20952_26 : GEN_1469;
  assign GEN_1471 = 9'h1b == T_24222 ? T_20952_27 : GEN_1470;
  assign GEN_1472 = 9'h1c == T_24222 ? T_20952_28 : GEN_1471;
  assign GEN_1473 = 9'h1d == T_24222 ? T_20952_29 : GEN_1472;
  assign GEN_1474 = 9'h1e == T_24222 ? T_20952_30 : GEN_1473;
  assign GEN_1475 = 9'h1f == T_24222 ? T_20952_31 : GEN_1474;
  assign GEN_1476 = 9'h20 == T_24222 ? T_20952_32 : GEN_1475;
  assign GEN_1477 = 9'h21 == T_24222 ? T_20952_33 : GEN_1476;
  assign GEN_1478 = 9'h22 == T_24222 ? T_20952_34 : GEN_1477;
  assign GEN_1479 = 9'h23 == T_24222 ? T_20952_35 : GEN_1478;
  assign GEN_1480 = 9'h24 == T_24222 ? T_20952_36 : GEN_1479;
  assign GEN_1481 = 9'h25 == T_24222 ? T_20952_37 : GEN_1480;
  assign GEN_1482 = 9'h26 == T_24222 ? T_20952_38 : GEN_1481;
  assign GEN_1483 = 9'h27 == T_24222 ? T_20952_39 : GEN_1482;
  assign GEN_1484 = 9'h28 == T_24222 ? T_20952_40 : GEN_1483;
  assign GEN_1485 = 9'h29 == T_24222 ? T_20952_41 : GEN_1484;
  assign GEN_1486 = 9'h2a == T_24222 ? T_20952_42 : GEN_1485;
  assign GEN_1487 = 9'h2b == T_24222 ? T_20952_43 : GEN_1486;
  assign GEN_1488 = 9'h2c == T_24222 ? T_20952_44 : GEN_1487;
  assign GEN_1489 = 9'h2d == T_24222 ? T_20952_45 : GEN_1488;
  assign GEN_1490 = 9'h2e == T_24222 ? T_20952_46 : GEN_1489;
  assign GEN_1491 = 9'h2f == T_24222 ? T_20952_47 : GEN_1490;
  assign GEN_1492 = 9'h30 == T_24222 ? T_20952_48 : GEN_1491;
  assign GEN_1493 = 9'h31 == T_24222 ? T_20952_49 : GEN_1492;
  assign GEN_1494 = 9'h32 == T_24222 ? T_20952_50 : GEN_1493;
  assign GEN_1495 = 9'h33 == T_24222 ? T_20952_51 : GEN_1494;
  assign GEN_1496 = 9'h34 == T_24222 ? T_20952_52 : GEN_1495;
  assign GEN_1497 = 9'h35 == T_24222 ? T_20952_53 : GEN_1496;
  assign GEN_1498 = 9'h36 == T_24222 ? T_20952_54 : GEN_1497;
  assign GEN_1499 = 9'h37 == T_24222 ? T_20952_55 : GEN_1498;
  assign GEN_1500 = 9'h38 == T_24222 ? T_20952_56 : GEN_1499;
  assign GEN_1501 = 9'h39 == T_24222 ? T_20952_57 : GEN_1500;
  assign GEN_1502 = 9'h3a == T_24222 ? T_20952_58 : GEN_1501;
  assign GEN_1503 = 9'h3b == T_24222 ? T_20952_59 : GEN_1502;
  assign GEN_1504 = 9'h3c == T_24222 ? T_20952_60 : GEN_1503;
  assign GEN_1505 = 9'h3d == T_24222 ? T_20952_61 : GEN_1504;
  assign GEN_1506 = 9'h3e == T_24222 ? T_20952_62 : GEN_1505;
  assign GEN_1507 = 9'h3f == T_24222 ? T_20952_63 : GEN_1506;
  assign GEN_1508 = 9'h40 == T_24222 ? T_20952_64 : GEN_1507;
  assign GEN_1509 = 9'h41 == T_24222 ? T_20952_65 : GEN_1508;
  assign GEN_1510 = 9'h42 == T_24222 ? T_20952_66 : GEN_1509;
  assign GEN_1511 = 9'h43 == T_24222 ? T_20952_67 : GEN_1510;
  assign GEN_1512 = 9'h44 == T_24222 ? T_20952_68 : GEN_1511;
  assign GEN_1513 = 9'h45 == T_24222 ? T_20952_69 : GEN_1512;
  assign GEN_1514 = 9'h46 == T_24222 ? T_20952_70 : GEN_1513;
  assign GEN_1515 = 9'h47 == T_24222 ? T_20952_71 : GEN_1514;
  assign GEN_1516 = 9'h48 == T_24222 ? T_20952_72 : GEN_1515;
  assign GEN_1517 = 9'h49 == T_24222 ? T_20952_73 : GEN_1516;
  assign GEN_1518 = 9'h4a == T_24222 ? T_20952_74 : GEN_1517;
  assign GEN_1519 = 9'h4b == T_24222 ? T_20952_75 : GEN_1518;
  assign GEN_1520 = 9'h4c == T_24222 ? T_20952_76 : GEN_1519;
  assign GEN_1521 = 9'h4d == T_24222 ? T_20952_77 : GEN_1520;
  assign GEN_1522 = 9'h4e == T_24222 ? T_20952_78 : GEN_1521;
  assign GEN_1523 = 9'h4f == T_24222 ? T_20952_79 : GEN_1522;
  assign GEN_1524 = 9'h50 == T_24222 ? T_20952_80 : GEN_1523;
  assign GEN_1525 = 9'h51 == T_24222 ? T_20952_81 : GEN_1524;
  assign GEN_1526 = 9'h52 == T_24222 ? T_20952_82 : GEN_1525;
  assign GEN_1527 = 9'h53 == T_24222 ? T_20952_83 : GEN_1526;
  assign GEN_1528 = 9'h54 == T_24222 ? T_20952_84 : GEN_1527;
  assign GEN_1529 = 9'h55 == T_24222 ? T_20952_85 : GEN_1528;
  assign GEN_1530 = 9'h56 == T_24222 ? T_20952_86 : GEN_1529;
  assign GEN_1531 = 9'h57 == T_24222 ? T_20952_87 : GEN_1530;
  assign GEN_1532 = 9'h58 == T_24222 ? T_20952_88 : GEN_1531;
  assign GEN_1533 = 9'h59 == T_24222 ? T_20952_89 : GEN_1532;
  assign GEN_1534 = 9'h5a == T_24222 ? T_20952_90 : GEN_1533;
  assign GEN_1535 = 9'h5b == T_24222 ? T_20952_91 : GEN_1534;
  assign GEN_1536 = 9'h5c == T_24222 ? T_20952_92 : GEN_1535;
  assign GEN_1537 = 9'h5d == T_24222 ? T_20952_93 : GEN_1536;
  assign GEN_1538 = 9'h5e == T_24222 ? T_20952_94 : GEN_1537;
  assign GEN_1539 = 9'h5f == T_24222 ? T_20952_95 : GEN_1538;
  assign GEN_1540 = 9'h60 == T_24222 ? T_20952_96 : GEN_1539;
  assign GEN_1541 = 9'h61 == T_24222 ? T_20952_97 : GEN_1540;
  assign GEN_1542 = 9'h62 == T_24222 ? T_20952_98 : GEN_1541;
  assign GEN_1543 = 9'h63 == T_24222 ? T_20952_99 : GEN_1542;
  assign GEN_1544 = 9'h64 == T_24222 ? T_20952_100 : GEN_1543;
  assign GEN_1545 = 9'h65 == T_24222 ? T_20952_101 : GEN_1544;
  assign GEN_1546 = 9'h66 == T_24222 ? T_20952_102 : GEN_1545;
  assign GEN_1547 = 9'h67 == T_24222 ? T_20952_103 : GEN_1546;
  assign GEN_1548 = 9'h68 == T_24222 ? T_20952_104 : GEN_1547;
  assign GEN_1549 = 9'h69 == T_24222 ? T_20952_105 : GEN_1548;
  assign GEN_1550 = 9'h6a == T_24222 ? T_20952_106 : GEN_1549;
  assign GEN_1551 = 9'h6b == T_24222 ? T_20952_107 : GEN_1550;
  assign GEN_1552 = 9'h6c == T_24222 ? T_20952_108 : GEN_1551;
  assign GEN_1553 = 9'h6d == T_24222 ? T_20952_109 : GEN_1552;
  assign GEN_1554 = 9'h6e == T_24222 ? T_20952_110 : GEN_1553;
  assign GEN_1555 = 9'h6f == T_24222 ? T_20952_111 : GEN_1554;
  assign GEN_1556 = 9'h70 == T_24222 ? T_20952_112 : GEN_1555;
  assign GEN_1557 = 9'h71 == T_24222 ? T_20952_113 : GEN_1556;
  assign GEN_1558 = 9'h72 == T_24222 ? T_20952_114 : GEN_1557;
  assign GEN_1559 = 9'h73 == T_24222 ? T_20952_115 : GEN_1558;
  assign GEN_1560 = 9'h74 == T_24222 ? T_20952_116 : GEN_1559;
  assign GEN_1561 = 9'h75 == T_24222 ? T_20952_117 : GEN_1560;
  assign GEN_1562 = 9'h76 == T_24222 ? T_20952_118 : GEN_1561;
  assign GEN_1563 = 9'h77 == T_24222 ? T_20952_119 : GEN_1562;
  assign GEN_1564 = 9'h78 == T_24222 ? T_20952_120 : GEN_1563;
  assign GEN_1565 = 9'h79 == T_24222 ? T_20952_121 : GEN_1564;
  assign GEN_1566 = 9'h7a == T_24222 ? T_20952_122 : GEN_1565;
  assign GEN_1567 = 9'h7b == T_24222 ? T_20952_123 : GEN_1566;
  assign GEN_1568 = 9'h7c == T_24222 ? T_20952_124 : GEN_1567;
  assign GEN_1569 = 9'h7d == T_24222 ? T_20952_125 : GEN_1568;
  assign GEN_1570 = 9'h7e == T_24222 ? T_20952_126 : GEN_1569;
  assign GEN_1571 = 9'h7f == T_24222 ? T_20952_127 : GEN_1570;
  assign GEN_1572 = 9'h80 == T_24222 ? T_20952_128 : GEN_1571;
  assign GEN_1573 = 9'h81 == T_24222 ? T_20952_129 : GEN_1572;
  assign GEN_1574 = 9'h82 == T_24222 ? T_20952_130 : GEN_1573;
  assign GEN_1575 = 9'h83 == T_24222 ? T_20952_131 : GEN_1574;
  assign GEN_1576 = 9'h84 == T_24222 ? T_20952_132 : GEN_1575;
  assign GEN_1577 = 9'h85 == T_24222 ? T_20952_133 : GEN_1576;
  assign GEN_1578 = 9'h86 == T_24222 ? T_20952_134 : GEN_1577;
  assign GEN_1579 = 9'h87 == T_24222 ? T_20952_135 : GEN_1578;
  assign GEN_1580 = 9'h88 == T_24222 ? T_20952_136 : GEN_1579;
  assign GEN_1581 = 9'h89 == T_24222 ? T_20952_137 : GEN_1580;
  assign GEN_1582 = 9'h8a == T_24222 ? T_20952_138 : GEN_1581;
  assign GEN_1583 = 9'h8b == T_24222 ? T_20952_139 : GEN_1582;
  assign GEN_1584 = 9'h8c == T_24222 ? T_20952_140 : GEN_1583;
  assign GEN_1585 = 9'h8d == T_24222 ? T_20952_141 : GEN_1584;
  assign GEN_1586 = 9'h8e == T_24222 ? T_20952_142 : GEN_1585;
  assign GEN_1587 = 9'h8f == T_24222 ? T_20952_143 : GEN_1586;
  assign GEN_1588 = 9'h90 == T_24222 ? T_20952_144 : GEN_1587;
  assign GEN_1589 = 9'h91 == T_24222 ? T_20952_145 : GEN_1588;
  assign GEN_1590 = 9'h92 == T_24222 ? T_20952_146 : GEN_1589;
  assign GEN_1591 = 9'h93 == T_24222 ? T_20952_147 : GEN_1590;
  assign GEN_1592 = 9'h94 == T_24222 ? T_20952_148 : GEN_1591;
  assign GEN_1593 = 9'h95 == T_24222 ? T_20952_149 : GEN_1592;
  assign GEN_1594 = 9'h96 == T_24222 ? T_20952_150 : GEN_1593;
  assign GEN_1595 = 9'h97 == T_24222 ? T_20952_151 : GEN_1594;
  assign GEN_1596 = 9'h98 == T_24222 ? T_20952_152 : GEN_1595;
  assign GEN_1597 = 9'h99 == T_24222 ? T_20952_153 : GEN_1596;
  assign GEN_1598 = 9'h9a == T_24222 ? T_20952_154 : GEN_1597;
  assign GEN_1599 = 9'h9b == T_24222 ? T_20952_155 : GEN_1598;
  assign GEN_1600 = 9'h9c == T_24222 ? T_20952_156 : GEN_1599;
  assign GEN_1601 = 9'h9d == T_24222 ? T_20952_157 : GEN_1600;
  assign GEN_1602 = 9'h9e == T_24222 ? T_20952_158 : GEN_1601;
  assign GEN_1603 = 9'h9f == T_24222 ? T_20952_159 : GEN_1602;
  assign GEN_1604 = 9'ha0 == T_24222 ? T_20952_160 : GEN_1603;
  assign GEN_1605 = 9'ha1 == T_24222 ? T_20952_161 : GEN_1604;
  assign GEN_1606 = 9'ha2 == T_24222 ? T_20952_162 : GEN_1605;
  assign GEN_1607 = 9'ha3 == T_24222 ? T_20952_163 : GEN_1606;
  assign GEN_1608 = 9'ha4 == T_24222 ? T_20952_164 : GEN_1607;
  assign GEN_1609 = 9'ha5 == T_24222 ? T_20952_165 : GEN_1608;
  assign GEN_1610 = 9'ha6 == T_24222 ? T_20952_166 : GEN_1609;
  assign GEN_1611 = 9'ha7 == T_24222 ? T_20952_167 : GEN_1610;
  assign GEN_1612 = 9'ha8 == T_24222 ? T_20952_168 : GEN_1611;
  assign GEN_1613 = 9'ha9 == T_24222 ? T_20952_169 : GEN_1612;
  assign GEN_1614 = 9'haa == T_24222 ? T_20952_170 : GEN_1613;
  assign GEN_1615 = 9'hab == T_24222 ? T_20952_171 : GEN_1614;
  assign GEN_1616 = 9'hac == T_24222 ? T_20952_172 : GEN_1615;
  assign GEN_1617 = 9'had == T_24222 ? T_20952_173 : GEN_1616;
  assign GEN_1618 = 9'hae == T_24222 ? T_20952_174 : GEN_1617;
  assign GEN_1619 = 9'haf == T_24222 ? T_20952_175 : GEN_1618;
  assign GEN_1620 = 9'hb0 == T_24222 ? T_20952_176 : GEN_1619;
  assign GEN_1621 = 9'hb1 == T_24222 ? T_20952_177 : GEN_1620;
  assign GEN_1622 = 9'hb2 == T_24222 ? T_20952_178 : GEN_1621;
  assign GEN_1623 = 9'hb3 == T_24222 ? T_20952_179 : GEN_1622;
  assign GEN_1624 = 9'hb4 == T_24222 ? T_20952_180 : GEN_1623;
  assign GEN_1625 = 9'hb5 == T_24222 ? T_20952_181 : GEN_1624;
  assign GEN_1626 = 9'hb6 == T_24222 ? T_20952_182 : GEN_1625;
  assign GEN_1627 = 9'hb7 == T_24222 ? T_20952_183 : GEN_1626;
  assign GEN_1628 = 9'hb8 == T_24222 ? T_20952_184 : GEN_1627;
  assign GEN_1629 = 9'hb9 == T_24222 ? T_20952_185 : GEN_1628;
  assign GEN_1630 = 9'hba == T_24222 ? T_20952_186 : GEN_1629;
  assign GEN_1631 = 9'hbb == T_24222 ? T_20952_187 : GEN_1630;
  assign GEN_1632 = 9'hbc == T_24222 ? T_20952_188 : GEN_1631;
  assign GEN_1633 = 9'hbd == T_24222 ? T_20952_189 : GEN_1632;
  assign GEN_1634 = 9'hbe == T_24222 ? T_20952_190 : GEN_1633;
  assign GEN_1635 = 9'hbf == T_24222 ? T_20952_191 : GEN_1634;
  assign GEN_1636 = 9'hc0 == T_24222 ? T_20952_192 : GEN_1635;
  assign GEN_1637 = 9'hc1 == T_24222 ? T_20952_193 : GEN_1636;
  assign GEN_1638 = 9'hc2 == T_24222 ? T_20952_194 : GEN_1637;
  assign GEN_1639 = 9'hc3 == T_24222 ? T_20952_195 : GEN_1638;
  assign GEN_1640 = 9'hc4 == T_24222 ? T_20952_196 : GEN_1639;
  assign GEN_1641 = 9'hc5 == T_24222 ? T_20952_197 : GEN_1640;
  assign GEN_1642 = 9'hc6 == T_24222 ? T_20952_198 : GEN_1641;
  assign GEN_1643 = 9'hc7 == T_24222 ? T_20952_199 : GEN_1642;
  assign GEN_1644 = 9'hc8 == T_24222 ? T_20952_200 : GEN_1643;
  assign GEN_1645 = 9'hc9 == T_24222 ? T_20952_201 : GEN_1644;
  assign GEN_1646 = 9'hca == T_24222 ? T_20952_202 : GEN_1645;
  assign GEN_1647 = 9'hcb == T_24222 ? T_20952_203 : GEN_1646;
  assign GEN_1648 = 9'hcc == T_24222 ? T_20952_204 : GEN_1647;
  assign GEN_1649 = 9'hcd == T_24222 ? T_20952_205 : GEN_1648;
  assign GEN_1650 = 9'hce == T_24222 ? T_20952_206 : GEN_1649;
  assign GEN_1651 = 9'hcf == T_24222 ? T_20952_207 : GEN_1650;
  assign GEN_1652 = 9'hd0 == T_24222 ? T_20952_208 : GEN_1651;
  assign GEN_1653 = 9'hd1 == T_24222 ? T_20952_209 : GEN_1652;
  assign GEN_1654 = 9'hd2 == T_24222 ? T_20952_210 : GEN_1653;
  assign GEN_1655 = 9'hd3 == T_24222 ? T_20952_211 : GEN_1654;
  assign GEN_1656 = 9'hd4 == T_24222 ? T_20952_212 : GEN_1655;
  assign GEN_1657 = 9'hd5 == T_24222 ? T_20952_213 : GEN_1656;
  assign GEN_1658 = 9'hd6 == T_24222 ? T_20952_214 : GEN_1657;
  assign GEN_1659 = 9'hd7 == T_24222 ? T_20952_215 : GEN_1658;
  assign GEN_1660 = 9'hd8 == T_24222 ? T_20952_216 : GEN_1659;
  assign GEN_1661 = 9'hd9 == T_24222 ? T_20952_217 : GEN_1660;
  assign GEN_1662 = 9'hda == T_24222 ? T_20952_218 : GEN_1661;
  assign GEN_1663 = 9'hdb == T_24222 ? T_20952_219 : GEN_1662;
  assign GEN_1664 = 9'hdc == T_24222 ? T_20952_220 : GEN_1663;
  assign GEN_1665 = 9'hdd == T_24222 ? T_20952_221 : GEN_1664;
  assign GEN_1666 = 9'hde == T_24222 ? T_20952_222 : GEN_1665;
  assign GEN_1667 = 9'hdf == T_24222 ? T_20952_223 : GEN_1666;
  assign GEN_1668 = 9'he0 == T_24222 ? T_20952_224 : GEN_1667;
  assign GEN_1669 = 9'he1 == T_24222 ? T_20952_225 : GEN_1668;
  assign GEN_1670 = 9'he2 == T_24222 ? T_20952_226 : GEN_1669;
  assign GEN_1671 = 9'he3 == T_24222 ? T_20952_227 : GEN_1670;
  assign GEN_1672 = 9'he4 == T_24222 ? T_20952_228 : GEN_1671;
  assign GEN_1673 = 9'he5 == T_24222 ? T_20952_229 : GEN_1672;
  assign GEN_1674 = 9'he6 == T_24222 ? T_20952_230 : GEN_1673;
  assign GEN_1675 = 9'he7 == T_24222 ? T_20952_231 : GEN_1674;
  assign GEN_1676 = 9'he8 == T_24222 ? T_20952_232 : GEN_1675;
  assign GEN_1677 = 9'he9 == T_24222 ? T_20952_233 : GEN_1676;
  assign GEN_1678 = 9'hea == T_24222 ? T_20952_234 : GEN_1677;
  assign GEN_1679 = 9'heb == T_24222 ? T_20952_235 : GEN_1678;
  assign GEN_1680 = 9'hec == T_24222 ? T_20952_236 : GEN_1679;
  assign GEN_1681 = 9'hed == T_24222 ? T_20952_237 : GEN_1680;
  assign GEN_1682 = 9'hee == T_24222 ? T_20952_238 : GEN_1681;
  assign GEN_1683 = 9'hef == T_24222 ? T_20952_239 : GEN_1682;
  assign GEN_1684 = 9'hf0 == T_24222 ? T_20952_240 : GEN_1683;
  assign GEN_1685 = 9'hf1 == T_24222 ? T_20952_241 : GEN_1684;
  assign GEN_1686 = 9'hf2 == T_24222 ? T_20952_242 : GEN_1685;
  assign GEN_1687 = 9'hf3 == T_24222 ? T_20952_243 : GEN_1686;
  assign GEN_1688 = 9'hf4 == T_24222 ? T_20952_244 : GEN_1687;
  assign GEN_1689 = 9'hf5 == T_24222 ? T_20952_245 : GEN_1688;
  assign GEN_1690 = 9'hf6 == T_24222 ? T_20952_246 : GEN_1689;
  assign GEN_1691 = 9'hf7 == T_24222 ? T_20952_247 : GEN_1690;
  assign GEN_1692 = 9'hf8 == T_24222 ? T_20952_248 : GEN_1691;
  assign GEN_1693 = 9'hf9 == T_24222 ? T_20952_249 : GEN_1692;
  assign GEN_1694 = 9'hfa == T_24222 ? T_20952_250 : GEN_1693;
  assign GEN_1695 = 9'hfb == T_24222 ? T_20952_251 : GEN_1694;
  assign GEN_1696 = 9'hfc == T_24222 ? T_20952_252 : GEN_1695;
  assign GEN_1697 = 9'hfd == T_24222 ? T_20952_253 : GEN_1696;
  assign GEN_1698 = 9'hfe == T_24222 ? T_20952_254 : GEN_1697;
  assign GEN_1699 = 9'hff == T_24222 ? T_20952_255 : GEN_1698;
  assign GEN_1700 = 9'h100 == T_24222 ? T_20952_256 : GEN_1699;
  assign GEN_1701 = 9'h101 == T_24222 ? T_20952_257 : GEN_1700;
  assign GEN_1702 = 9'h102 == T_24222 ? T_20952_258 : GEN_1701;
  assign GEN_1703 = 9'h103 == T_24222 ? T_20952_259 : GEN_1702;
  assign GEN_1704 = 9'h104 == T_24222 ? T_20952_260 : GEN_1703;
  assign GEN_1705 = 9'h105 == T_24222 ? T_20952_261 : GEN_1704;
  assign GEN_1706 = 9'h106 == T_24222 ? T_20952_262 : GEN_1705;
  assign GEN_1707 = 9'h107 == T_24222 ? T_20952_263 : GEN_1706;
  assign GEN_1708 = 9'h108 == T_24222 ? T_20952_264 : GEN_1707;
  assign GEN_1709 = 9'h109 == T_24222 ? T_20952_265 : GEN_1708;
  assign GEN_1710 = 9'h10a == T_24222 ? T_20952_266 : GEN_1709;
  assign GEN_1711 = 9'h10b == T_24222 ? T_20952_267 : GEN_1710;
  assign GEN_1712 = 9'h10c == T_24222 ? T_20952_268 : GEN_1711;
  assign GEN_1713 = 9'h10d == T_24222 ? T_20952_269 : GEN_1712;
  assign GEN_1714 = 9'h10e == T_24222 ? T_20952_270 : GEN_1713;
  assign GEN_1715 = 9'h10f == T_24222 ? T_20952_271 : GEN_1714;
  assign GEN_1716 = 9'h110 == T_24222 ? T_20952_272 : GEN_1715;
  assign GEN_1717 = 9'h111 == T_24222 ? T_20952_273 : GEN_1716;
  assign GEN_1718 = 9'h112 == T_24222 ? T_20952_274 : GEN_1717;
  assign GEN_1719 = 9'h113 == T_24222 ? T_20952_275 : GEN_1718;
  assign GEN_1720 = 9'h114 == T_24222 ? T_20952_276 : GEN_1719;
  assign GEN_1721 = 9'h115 == T_24222 ? T_20952_277 : GEN_1720;
  assign GEN_1722 = 9'h116 == T_24222 ? T_20952_278 : GEN_1721;
  assign GEN_1723 = 9'h117 == T_24222 ? T_20952_279 : GEN_1722;
  assign GEN_1724 = 9'h118 == T_24222 ? T_20952_280 : GEN_1723;
  assign GEN_1725 = 9'h119 == T_24222 ? T_20952_281 : GEN_1724;
  assign GEN_1726 = 9'h11a == T_24222 ? T_20952_282 : GEN_1725;
  assign GEN_1727 = 9'h11b == T_24222 ? T_20952_283 : GEN_1726;
  assign GEN_1728 = 9'h11c == T_24222 ? T_20952_284 : GEN_1727;
  assign GEN_1729 = 9'h11d == T_24222 ? T_20952_285 : GEN_1728;
  assign GEN_1730 = 9'h11e == T_24222 ? T_20952_286 : GEN_1729;
  assign GEN_1731 = 9'h11f == T_24222 ? T_20952_287 : GEN_1730;
  assign GEN_1732 = 9'h120 == T_24222 ? T_20952_288 : GEN_1731;
  assign GEN_1733 = 9'h121 == T_24222 ? T_20952_289 : GEN_1732;
  assign GEN_1734 = 9'h122 == T_24222 ? T_20952_290 : GEN_1733;
  assign GEN_1735 = 9'h123 == T_24222 ? T_20952_291 : GEN_1734;
  assign GEN_1736 = 9'h124 == T_24222 ? T_20952_292 : GEN_1735;
  assign GEN_1737 = 9'h125 == T_24222 ? T_20952_293 : GEN_1736;
  assign GEN_1738 = 9'h126 == T_24222 ? T_20952_294 : GEN_1737;
  assign GEN_1739 = 9'h127 == T_24222 ? T_20952_295 : GEN_1738;
  assign GEN_1740 = 9'h128 == T_24222 ? T_20952_296 : GEN_1739;
  assign GEN_1741 = 9'h129 == T_24222 ? T_20952_297 : GEN_1740;
  assign GEN_1742 = 9'h12a == T_24222 ? T_20952_298 : GEN_1741;
  assign GEN_1743 = 9'h12b == T_24222 ? T_20952_299 : GEN_1742;
  assign GEN_1744 = 9'h12c == T_24222 ? T_20952_300 : GEN_1743;
  assign GEN_1745 = 9'h12d == T_24222 ? T_20952_301 : GEN_1744;
  assign GEN_1746 = 9'h12e == T_24222 ? T_20952_302 : GEN_1745;
  assign GEN_1747 = 9'h12f == T_24222 ? T_20952_303 : GEN_1746;
  assign GEN_1748 = 9'h130 == T_24222 ? T_20952_304 : GEN_1747;
  assign GEN_1749 = 9'h131 == T_24222 ? T_20952_305 : GEN_1748;
  assign GEN_1750 = 9'h132 == T_24222 ? T_20952_306 : GEN_1749;
  assign GEN_1751 = 9'h133 == T_24222 ? T_20952_307 : GEN_1750;
  assign GEN_1752 = 9'h134 == T_24222 ? T_20952_308 : GEN_1751;
  assign GEN_1753 = 9'h135 == T_24222 ? T_20952_309 : GEN_1752;
  assign GEN_1754 = 9'h136 == T_24222 ? T_20952_310 : GEN_1753;
  assign GEN_1755 = 9'h137 == T_24222 ? T_20952_311 : GEN_1754;
  assign GEN_1756 = 9'h138 == T_24222 ? T_20952_312 : GEN_1755;
  assign GEN_1757 = 9'h139 == T_24222 ? T_20952_313 : GEN_1756;
  assign GEN_1758 = 9'h13a == T_24222 ? T_20952_314 : GEN_1757;
  assign GEN_1759 = 9'h13b == T_24222 ? T_20952_315 : GEN_1758;
  assign GEN_1760 = 9'h13c == T_24222 ? T_20952_316 : GEN_1759;
  assign GEN_1761 = 9'h13d == T_24222 ? T_20952_317 : GEN_1760;
  assign GEN_1762 = 9'h13e == T_24222 ? T_20952_318 : GEN_1761;
  assign GEN_1763 = 9'h13f == T_24222 ? T_20952_319 : GEN_1762;
  assign GEN_1764 = 9'h140 == T_24222 ? T_20952_320 : GEN_1763;
  assign GEN_1765 = 9'h141 == T_24222 ? T_20952_321 : GEN_1764;
  assign GEN_1766 = 9'h142 == T_24222 ? T_20952_322 : GEN_1765;
  assign GEN_1767 = 9'h143 == T_24222 ? T_20952_323 : GEN_1766;
  assign GEN_1768 = 9'h144 == T_24222 ? T_20952_324 : GEN_1767;
  assign GEN_1769 = 9'h145 == T_24222 ? T_20952_325 : GEN_1768;
  assign GEN_1770 = 9'h146 == T_24222 ? T_20952_326 : GEN_1769;
  assign GEN_1771 = 9'h147 == T_24222 ? T_20952_327 : GEN_1770;
  assign GEN_1772 = 9'h148 == T_24222 ? T_20952_328 : GEN_1771;
  assign GEN_1773 = 9'h149 == T_24222 ? T_20952_329 : GEN_1772;
  assign GEN_1774 = 9'h14a == T_24222 ? T_20952_330 : GEN_1773;
  assign GEN_1775 = 9'h14b == T_24222 ? T_20952_331 : GEN_1774;
  assign GEN_1776 = 9'h14c == T_24222 ? T_20952_332 : GEN_1775;
  assign GEN_1777 = 9'h14d == T_24222 ? T_20952_333 : GEN_1776;
  assign GEN_1778 = 9'h14e == T_24222 ? T_20952_334 : GEN_1777;
  assign GEN_1779 = 9'h14f == T_24222 ? T_20952_335 : GEN_1778;
  assign GEN_1780 = 9'h150 == T_24222 ? T_20952_336 : GEN_1779;
  assign GEN_1781 = 9'h151 == T_24222 ? T_20952_337 : GEN_1780;
  assign GEN_1782 = 9'h152 == T_24222 ? T_20952_338 : GEN_1781;
  assign GEN_1783 = 9'h153 == T_24222 ? T_20952_339 : GEN_1782;
  assign GEN_1784 = 9'h154 == T_24222 ? T_20952_340 : GEN_1783;
  assign GEN_1785 = 9'h155 == T_24222 ? T_20952_341 : GEN_1784;
  assign GEN_1786 = 9'h156 == T_24222 ? T_20952_342 : GEN_1785;
  assign GEN_1787 = 9'h157 == T_24222 ? T_20952_343 : GEN_1786;
  assign GEN_1788 = 9'h158 == T_24222 ? T_20952_344 : GEN_1787;
  assign GEN_1789 = 9'h159 == T_24222 ? T_20952_345 : GEN_1788;
  assign GEN_1790 = 9'h15a == T_24222 ? T_20952_346 : GEN_1789;
  assign GEN_1791 = 9'h15b == T_24222 ? T_20952_347 : GEN_1790;
  assign GEN_1792 = 9'h15c == T_24222 ? T_20952_348 : GEN_1791;
  assign GEN_1793 = 9'h15d == T_24222 ? T_20952_349 : GEN_1792;
  assign GEN_1794 = 9'h15e == T_24222 ? T_20952_350 : GEN_1793;
  assign GEN_1795 = 9'h15f == T_24222 ? T_20952_351 : GEN_1794;
  assign GEN_1796 = 9'h160 == T_24222 ? T_20952_352 : GEN_1795;
  assign GEN_1797 = 9'h161 == T_24222 ? T_20952_353 : GEN_1796;
  assign GEN_1798 = 9'h162 == T_24222 ? T_20952_354 : GEN_1797;
  assign GEN_1799 = 9'h163 == T_24222 ? T_20952_355 : GEN_1798;
  assign GEN_1800 = 9'h164 == T_24222 ? T_20952_356 : GEN_1799;
  assign GEN_1801 = 9'h165 == T_24222 ? T_20952_357 : GEN_1800;
  assign GEN_1802 = 9'h166 == T_24222 ? T_20952_358 : GEN_1801;
  assign GEN_1803 = 9'h167 == T_24222 ? T_20952_359 : GEN_1802;
  assign GEN_1804 = 9'h168 == T_24222 ? T_20952_360 : GEN_1803;
  assign GEN_1805 = 9'h169 == T_24222 ? T_20952_361 : GEN_1804;
  assign GEN_1806 = 9'h16a == T_24222 ? T_20952_362 : GEN_1805;
  assign GEN_1807 = 9'h16b == T_24222 ? T_20952_363 : GEN_1806;
  assign GEN_1808 = 9'h16c == T_24222 ? T_20952_364 : GEN_1807;
  assign GEN_1809 = 9'h16d == T_24222 ? T_20952_365 : GEN_1808;
  assign GEN_1810 = 9'h16e == T_24222 ? T_20952_366 : GEN_1809;
  assign GEN_1811 = 9'h16f == T_24222 ? T_20952_367 : GEN_1810;
  assign GEN_1812 = 9'h170 == T_24222 ? T_20952_368 : GEN_1811;
  assign GEN_1813 = 9'h171 == T_24222 ? T_20952_369 : GEN_1812;
  assign GEN_1814 = 9'h172 == T_24222 ? T_20952_370 : GEN_1813;
  assign GEN_1815 = 9'h173 == T_24222 ? T_20952_371 : GEN_1814;
  assign GEN_1816 = 9'h174 == T_24222 ? T_20952_372 : GEN_1815;
  assign GEN_1817 = 9'h175 == T_24222 ? T_20952_373 : GEN_1816;
  assign GEN_1818 = 9'h176 == T_24222 ? T_20952_374 : GEN_1817;
  assign GEN_1819 = 9'h177 == T_24222 ? T_20952_375 : GEN_1818;
  assign GEN_1820 = 9'h178 == T_24222 ? T_20952_376 : GEN_1819;
  assign GEN_1821 = 9'h179 == T_24222 ? T_20952_377 : GEN_1820;
  assign GEN_1822 = 9'h17a == T_24222 ? T_20952_378 : GEN_1821;
  assign GEN_1823 = 9'h17b == T_24222 ? T_20952_379 : GEN_1822;
  assign GEN_1824 = 9'h17c == T_24222 ? T_20952_380 : GEN_1823;
  assign GEN_1825 = 9'h17d == T_24222 ? T_20952_381 : GEN_1824;
  assign GEN_1826 = 9'h17e == T_24222 ? T_20952_382 : GEN_1825;
  assign GEN_1827 = 9'h17f == T_24222 ? T_20952_383 : GEN_1826;
  assign GEN_1828 = 9'h180 == T_24222 ? T_20952_384 : GEN_1827;
  assign GEN_1829 = 9'h181 == T_24222 ? T_20952_385 : GEN_1828;
  assign GEN_1830 = 9'h182 == T_24222 ? T_20952_386 : GEN_1829;
  assign GEN_1831 = 9'h183 == T_24222 ? T_20952_387 : GEN_1830;
  assign GEN_1832 = 9'h184 == T_24222 ? T_20952_388 : GEN_1831;
  assign GEN_1833 = 9'h185 == T_24222 ? T_20952_389 : GEN_1832;
  assign GEN_1834 = 9'h186 == T_24222 ? T_20952_390 : GEN_1833;
  assign GEN_1835 = 9'h187 == T_24222 ? T_20952_391 : GEN_1834;
  assign GEN_1836 = 9'h188 == T_24222 ? T_20952_392 : GEN_1835;
  assign GEN_1837 = 9'h189 == T_24222 ? T_20952_393 : GEN_1836;
  assign GEN_1838 = 9'h18a == T_24222 ? T_20952_394 : GEN_1837;
  assign GEN_1839 = 9'h18b == T_24222 ? T_20952_395 : GEN_1838;
  assign GEN_1840 = 9'h18c == T_24222 ? T_20952_396 : GEN_1839;
  assign GEN_1841 = 9'h18d == T_24222 ? T_20952_397 : GEN_1840;
  assign GEN_1842 = 9'h18e == T_24222 ? T_20952_398 : GEN_1841;
  assign GEN_1843 = 9'h18f == T_24222 ? T_20952_399 : GEN_1842;
  assign GEN_1844 = 9'h190 == T_24222 ? T_20952_400 : GEN_1843;
  assign GEN_1845 = 9'h191 == T_24222 ? T_20952_401 : GEN_1844;
  assign GEN_1846 = 9'h192 == T_24222 ? T_20952_402 : GEN_1845;
  assign GEN_1847 = 9'h193 == T_24222 ? T_20952_403 : GEN_1846;
  assign GEN_1848 = 9'h194 == T_24222 ? T_20952_404 : GEN_1847;
  assign GEN_1849 = 9'h195 == T_24222 ? T_20952_405 : GEN_1848;
  assign GEN_1850 = 9'h196 == T_24222 ? T_20952_406 : GEN_1849;
  assign GEN_1851 = 9'h197 == T_24222 ? T_20952_407 : GEN_1850;
  assign GEN_1852 = 9'h198 == T_24222 ? T_20952_408 : GEN_1851;
  assign GEN_1853 = 9'h199 == T_24222 ? T_20952_409 : GEN_1852;
  assign GEN_1854 = 9'h19a == T_24222 ? T_20952_410 : GEN_1853;
  assign GEN_1855 = 9'h19b == T_24222 ? T_20952_411 : GEN_1854;
  assign GEN_1856 = 9'h19c == T_24222 ? T_20952_412 : GEN_1855;
  assign GEN_1857 = 9'h19d == T_24222 ? T_20952_413 : GEN_1856;
  assign GEN_1858 = 9'h19e == T_24222 ? T_20952_414 : GEN_1857;
  assign GEN_1859 = 9'h19f == T_24222 ? T_20952_415 : GEN_1858;
  assign GEN_1860 = 9'h1a0 == T_24222 ? T_20952_416 : GEN_1859;
  assign GEN_1861 = 9'h1a1 == T_24222 ? T_20952_417 : GEN_1860;
  assign GEN_1862 = 9'h1a2 == T_24222 ? T_20952_418 : GEN_1861;
  assign GEN_1863 = 9'h1a3 == T_24222 ? T_20952_419 : GEN_1862;
  assign GEN_1864 = 9'h1a4 == T_24222 ? T_20952_420 : GEN_1863;
  assign GEN_1865 = 9'h1a5 == T_24222 ? T_20952_421 : GEN_1864;
  assign GEN_1866 = 9'h1a6 == T_24222 ? T_20952_422 : GEN_1865;
  assign GEN_1867 = 9'h1a7 == T_24222 ? T_20952_423 : GEN_1866;
  assign GEN_1868 = 9'h1a8 == T_24222 ? T_20952_424 : GEN_1867;
  assign GEN_1869 = 9'h1a9 == T_24222 ? T_20952_425 : GEN_1868;
  assign GEN_1870 = 9'h1aa == T_24222 ? T_20952_426 : GEN_1869;
  assign GEN_1871 = 9'h1ab == T_24222 ? T_20952_427 : GEN_1870;
  assign GEN_1872 = 9'h1ac == T_24222 ? T_20952_428 : GEN_1871;
  assign GEN_1873 = 9'h1ad == T_24222 ? T_20952_429 : GEN_1872;
  assign GEN_1874 = 9'h1ae == T_24222 ? T_20952_430 : GEN_1873;
  assign GEN_1875 = 9'h1af == T_24222 ? T_20952_431 : GEN_1874;
  assign GEN_1876 = 9'h1b0 == T_24222 ? T_20952_432 : GEN_1875;
  assign GEN_1877 = 9'h1b1 == T_24222 ? T_20952_433 : GEN_1876;
  assign GEN_1878 = 9'h1b2 == T_24222 ? T_20952_434 : GEN_1877;
  assign GEN_1879 = 9'h1b3 == T_24222 ? T_20952_435 : GEN_1878;
  assign GEN_1880 = 9'h1b4 == T_24222 ? T_20952_436 : GEN_1879;
  assign GEN_1881 = 9'h1b5 == T_24222 ? T_20952_437 : GEN_1880;
  assign GEN_1882 = 9'h1b6 == T_24222 ? T_20952_438 : GEN_1881;
  assign GEN_1883 = 9'h1b7 == T_24222 ? T_20952_439 : GEN_1882;
  assign GEN_1884 = 9'h1b8 == T_24222 ? T_20952_440 : GEN_1883;
  assign GEN_1885 = 9'h1b9 == T_24222 ? T_20952_441 : GEN_1884;
  assign GEN_1886 = 9'h1ba == T_24222 ? T_20952_442 : GEN_1885;
  assign GEN_1887 = 9'h1bb == T_24222 ? T_20952_443 : GEN_1886;
  assign GEN_1888 = 9'h1bc == T_24222 ? T_20952_444 : GEN_1887;
  assign GEN_1889 = 9'h1bd == T_24222 ? T_20952_445 : GEN_1888;
  assign GEN_1890 = 9'h1be == T_24222 ? T_20952_446 : GEN_1889;
  assign GEN_1891 = 9'h1bf == T_24222 ? T_20952_447 : GEN_1890;
  assign GEN_1892 = 9'h1c0 == T_24222 ? T_20952_448 : GEN_1891;
  assign GEN_1893 = 9'h1c1 == T_24222 ? T_20952_449 : GEN_1892;
  assign GEN_1894 = 9'h1c2 == T_24222 ? T_20952_450 : GEN_1893;
  assign GEN_1895 = 9'h1c3 == T_24222 ? T_20952_451 : GEN_1894;
  assign GEN_1896 = 9'h1c4 == T_24222 ? T_20952_452 : GEN_1895;
  assign GEN_1897 = 9'h1c5 == T_24222 ? T_20952_453 : GEN_1896;
  assign GEN_1898 = 9'h1c6 == T_24222 ? T_20952_454 : GEN_1897;
  assign GEN_1899 = 9'h1c7 == T_24222 ? T_20952_455 : GEN_1898;
  assign GEN_1900 = 9'h1c8 == T_24222 ? T_20952_456 : GEN_1899;
  assign GEN_1901 = 9'h1c9 == T_24222 ? T_20952_457 : GEN_1900;
  assign GEN_1902 = 9'h1ca == T_24222 ? T_20952_458 : GEN_1901;
  assign GEN_1903 = 9'h1cb == T_24222 ? T_20952_459 : GEN_1902;
  assign GEN_1904 = 9'h1cc == T_24222 ? T_20952_460 : GEN_1903;
  assign GEN_1905 = 9'h1cd == T_24222 ? T_20952_461 : GEN_1904;
  assign GEN_1906 = 9'h1ce == T_24222 ? T_20952_462 : GEN_1905;
  assign GEN_1907 = 9'h1cf == T_24222 ? T_20952_463 : GEN_1906;
  assign GEN_1908 = 9'h1d0 == T_24222 ? T_20952_464 : GEN_1907;
  assign GEN_1909 = 9'h1d1 == T_24222 ? T_20952_465 : GEN_1908;
  assign GEN_1910 = 9'h1d2 == T_24222 ? T_20952_466 : GEN_1909;
  assign GEN_1911 = 9'h1d3 == T_24222 ? T_20952_467 : GEN_1910;
  assign GEN_1912 = 9'h1d4 == T_24222 ? T_20952_468 : GEN_1911;
  assign GEN_1913 = 9'h1d5 == T_24222 ? T_20952_469 : GEN_1912;
  assign GEN_1914 = 9'h1d6 == T_24222 ? T_20952_470 : GEN_1913;
  assign GEN_1915 = 9'h1d7 == T_24222 ? T_20952_471 : GEN_1914;
  assign GEN_1916 = 9'h1d8 == T_24222 ? T_20952_472 : GEN_1915;
  assign GEN_1917 = 9'h1d9 == T_24222 ? T_20952_473 : GEN_1916;
  assign GEN_1918 = 9'h1da == T_24222 ? T_20952_474 : GEN_1917;
  assign GEN_1919 = 9'h1db == T_24222 ? T_20952_475 : GEN_1918;
  assign GEN_1920 = 9'h1dc == T_24222 ? T_20952_476 : GEN_1919;
  assign GEN_1921 = 9'h1dd == T_24222 ? T_20952_477 : GEN_1920;
  assign GEN_1922 = 9'h1de == T_24222 ? T_20952_478 : GEN_1921;
  assign GEN_1923 = 9'h1df == T_24222 ? T_20952_479 : GEN_1922;
  assign GEN_1924 = 9'h1e0 == T_24222 ? T_20952_480 : GEN_1923;
  assign GEN_1925 = 9'h1e1 == T_24222 ? T_20952_481 : GEN_1924;
  assign GEN_1926 = 9'h1e2 == T_24222 ? T_20952_482 : GEN_1925;
  assign GEN_1927 = 9'h1e3 == T_24222 ? T_20952_483 : GEN_1926;
  assign GEN_1928 = 9'h1e4 == T_24222 ? T_20952_484 : GEN_1927;
  assign GEN_1929 = 9'h1e5 == T_24222 ? T_20952_485 : GEN_1928;
  assign GEN_1930 = 9'h1e6 == T_24222 ? T_20952_486 : GEN_1929;
  assign GEN_1931 = 9'h1e7 == T_24222 ? T_20952_487 : GEN_1930;
  assign GEN_1932 = 9'h1e8 == T_24222 ? T_20952_488 : GEN_1931;
  assign GEN_1933 = 9'h1e9 == T_24222 ? T_20952_489 : GEN_1932;
  assign GEN_1934 = 9'h1ea == T_24222 ? T_20952_490 : GEN_1933;
  assign GEN_1935 = 9'h1eb == T_24222 ? T_20952_491 : GEN_1934;
  assign GEN_1936 = 9'h1ec == T_24222 ? T_20952_492 : GEN_1935;
  assign GEN_1937 = 9'h1ed == T_24222 ? T_20952_493 : GEN_1936;
  assign GEN_1938 = 9'h1ee == T_24222 ? T_20952_494 : GEN_1937;
  assign GEN_1939 = 9'h1ef == T_24222 ? T_20952_495 : GEN_1938;
  assign GEN_1940 = 9'h1f0 == T_24222 ? T_20952_496 : GEN_1939;
  assign GEN_1941 = 9'h1f1 == T_24222 ? T_20952_497 : GEN_1940;
  assign GEN_1942 = 9'h1f2 == T_24222 ? T_20952_498 : GEN_1941;
  assign GEN_1943 = 9'h1f3 == T_24222 ? T_20952_499 : GEN_1942;
  assign GEN_1944 = 9'h1f4 == T_24222 ? T_20952_500 : GEN_1943;
  assign GEN_1945 = 9'h1f5 == T_24222 ? T_20952_501 : GEN_1944;
  assign GEN_1946 = 9'h1f6 == T_24222 ? T_20952_502 : GEN_1945;
  assign GEN_1947 = 9'h1f7 == T_24222 ? T_20952_503 : GEN_1946;
  assign GEN_1948 = 9'h1f8 == T_24222 ? T_20952_504 : GEN_1947;
  assign GEN_1949 = 9'h1f9 == T_24222 ? T_20952_505 : GEN_1948;
  assign GEN_1950 = 9'h1fa == T_24222 ? T_20952_506 : GEN_1949;
  assign GEN_1951 = 9'h1fb == T_24222 ? T_20952_507 : GEN_1950;
  assign GEN_1952 = 9'h1fc == T_24222 ? T_20952_508 : GEN_1951;
  assign GEN_1953 = 9'h1fd == T_24222 ? T_20952_509 : GEN_1952;
  assign GEN_1954 = 9'h1fe == T_24222 ? T_20952_510 : GEN_1953;
  assign GEN_1955 = 9'h1ff == T_24222 ? T_20952_511 : GEN_1954;
  assign GEN_6 = GEN_2466;
  assign GEN_1956 = 9'h1 == T_24222 ? T_23676_1 : T_23676_0;
  assign GEN_1957 = 9'h2 == T_24222 ? T_23676_2 : GEN_1956;
  assign GEN_1958 = 9'h3 == T_24222 ? T_23676_3 : GEN_1957;
  assign GEN_1959 = 9'h4 == T_24222 ? T_23676_4 : GEN_1958;
  assign GEN_1960 = 9'h5 == T_24222 ? T_23676_5 : GEN_1959;
  assign GEN_1961 = 9'h6 == T_24222 ? T_23676_6 : GEN_1960;
  assign GEN_1962 = 9'h7 == T_24222 ? T_23676_7 : GEN_1961;
  assign GEN_1963 = 9'h8 == T_24222 ? T_23676_8 : GEN_1962;
  assign GEN_1964 = 9'h9 == T_24222 ? T_23676_9 : GEN_1963;
  assign GEN_1965 = 9'ha == T_24222 ? T_23676_10 : GEN_1964;
  assign GEN_1966 = 9'hb == T_24222 ? T_23676_11 : GEN_1965;
  assign GEN_1967 = 9'hc == T_24222 ? T_23676_12 : GEN_1966;
  assign GEN_1968 = 9'hd == T_24222 ? T_23676_13 : GEN_1967;
  assign GEN_1969 = 9'he == T_24222 ? T_23676_14 : GEN_1968;
  assign GEN_1970 = 9'hf == T_24222 ? T_23676_15 : GEN_1969;
  assign GEN_1971 = 9'h10 == T_24222 ? T_23676_16 : GEN_1970;
  assign GEN_1972 = 9'h11 == T_24222 ? T_23676_17 : GEN_1971;
  assign GEN_1973 = 9'h12 == T_24222 ? T_23676_18 : GEN_1972;
  assign GEN_1974 = 9'h13 == T_24222 ? T_23676_19 : GEN_1973;
  assign GEN_1975 = 9'h14 == T_24222 ? T_23676_20 : GEN_1974;
  assign GEN_1976 = 9'h15 == T_24222 ? T_23676_21 : GEN_1975;
  assign GEN_1977 = 9'h16 == T_24222 ? T_23676_22 : GEN_1976;
  assign GEN_1978 = 9'h17 == T_24222 ? T_23676_23 : GEN_1977;
  assign GEN_1979 = 9'h18 == T_24222 ? T_23676_24 : GEN_1978;
  assign GEN_1980 = 9'h19 == T_24222 ? T_23676_25 : GEN_1979;
  assign GEN_1981 = 9'h1a == T_24222 ? T_23676_26 : GEN_1980;
  assign GEN_1982 = 9'h1b == T_24222 ? T_23676_27 : GEN_1981;
  assign GEN_1983 = 9'h1c == T_24222 ? T_23676_28 : GEN_1982;
  assign GEN_1984 = 9'h1d == T_24222 ? T_23676_29 : GEN_1983;
  assign GEN_1985 = 9'h1e == T_24222 ? T_23676_30 : GEN_1984;
  assign GEN_1986 = 9'h1f == T_24222 ? T_23676_31 : GEN_1985;
  assign GEN_1987 = 9'h20 == T_24222 ? T_23676_32 : GEN_1986;
  assign GEN_1988 = 9'h21 == T_24222 ? T_23676_33 : GEN_1987;
  assign GEN_1989 = 9'h22 == T_24222 ? T_23676_34 : GEN_1988;
  assign GEN_1990 = 9'h23 == T_24222 ? T_23676_35 : GEN_1989;
  assign GEN_1991 = 9'h24 == T_24222 ? T_23676_36 : GEN_1990;
  assign GEN_1992 = 9'h25 == T_24222 ? T_23676_37 : GEN_1991;
  assign GEN_1993 = 9'h26 == T_24222 ? T_23676_38 : GEN_1992;
  assign GEN_1994 = 9'h27 == T_24222 ? T_23676_39 : GEN_1993;
  assign GEN_1995 = 9'h28 == T_24222 ? T_23676_40 : GEN_1994;
  assign GEN_1996 = 9'h29 == T_24222 ? T_23676_41 : GEN_1995;
  assign GEN_1997 = 9'h2a == T_24222 ? T_23676_42 : GEN_1996;
  assign GEN_1998 = 9'h2b == T_24222 ? T_23676_43 : GEN_1997;
  assign GEN_1999 = 9'h2c == T_24222 ? T_23676_44 : GEN_1998;
  assign GEN_2000 = 9'h2d == T_24222 ? T_23676_45 : GEN_1999;
  assign GEN_2001 = 9'h2e == T_24222 ? T_23676_46 : GEN_2000;
  assign GEN_2002 = 9'h2f == T_24222 ? T_23676_47 : GEN_2001;
  assign GEN_2003 = 9'h30 == T_24222 ? T_23676_48 : GEN_2002;
  assign GEN_2004 = 9'h31 == T_24222 ? T_23676_49 : GEN_2003;
  assign GEN_2005 = 9'h32 == T_24222 ? T_23676_50 : GEN_2004;
  assign GEN_2006 = 9'h33 == T_24222 ? T_23676_51 : GEN_2005;
  assign GEN_2007 = 9'h34 == T_24222 ? T_23676_52 : GEN_2006;
  assign GEN_2008 = 9'h35 == T_24222 ? T_23676_53 : GEN_2007;
  assign GEN_2009 = 9'h36 == T_24222 ? T_23676_54 : GEN_2008;
  assign GEN_2010 = 9'h37 == T_24222 ? T_23676_55 : GEN_2009;
  assign GEN_2011 = 9'h38 == T_24222 ? T_23676_56 : GEN_2010;
  assign GEN_2012 = 9'h39 == T_24222 ? T_23676_57 : GEN_2011;
  assign GEN_2013 = 9'h3a == T_24222 ? T_23676_58 : GEN_2012;
  assign GEN_2014 = 9'h3b == T_24222 ? T_23676_59 : GEN_2013;
  assign GEN_2015 = 9'h3c == T_24222 ? T_23676_60 : GEN_2014;
  assign GEN_2016 = 9'h3d == T_24222 ? T_23676_61 : GEN_2015;
  assign GEN_2017 = 9'h3e == T_24222 ? T_23676_62 : GEN_2016;
  assign GEN_2018 = 9'h3f == T_24222 ? T_23676_63 : GEN_2017;
  assign GEN_2019 = 9'h40 == T_24222 ? T_23676_64 : GEN_2018;
  assign GEN_2020 = 9'h41 == T_24222 ? T_23676_65 : GEN_2019;
  assign GEN_2021 = 9'h42 == T_24222 ? T_23676_66 : GEN_2020;
  assign GEN_2022 = 9'h43 == T_24222 ? T_23676_67 : GEN_2021;
  assign GEN_2023 = 9'h44 == T_24222 ? T_23676_68 : GEN_2022;
  assign GEN_2024 = 9'h45 == T_24222 ? T_23676_69 : GEN_2023;
  assign GEN_2025 = 9'h46 == T_24222 ? T_23676_70 : GEN_2024;
  assign GEN_2026 = 9'h47 == T_24222 ? T_23676_71 : GEN_2025;
  assign GEN_2027 = 9'h48 == T_24222 ? T_23676_72 : GEN_2026;
  assign GEN_2028 = 9'h49 == T_24222 ? T_23676_73 : GEN_2027;
  assign GEN_2029 = 9'h4a == T_24222 ? T_23676_74 : GEN_2028;
  assign GEN_2030 = 9'h4b == T_24222 ? T_23676_75 : GEN_2029;
  assign GEN_2031 = 9'h4c == T_24222 ? T_23676_76 : GEN_2030;
  assign GEN_2032 = 9'h4d == T_24222 ? T_23676_77 : GEN_2031;
  assign GEN_2033 = 9'h4e == T_24222 ? T_23676_78 : GEN_2032;
  assign GEN_2034 = 9'h4f == T_24222 ? T_23676_79 : GEN_2033;
  assign GEN_2035 = 9'h50 == T_24222 ? T_23676_80 : GEN_2034;
  assign GEN_2036 = 9'h51 == T_24222 ? T_23676_81 : GEN_2035;
  assign GEN_2037 = 9'h52 == T_24222 ? T_23676_82 : GEN_2036;
  assign GEN_2038 = 9'h53 == T_24222 ? T_23676_83 : GEN_2037;
  assign GEN_2039 = 9'h54 == T_24222 ? T_23676_84 : GEN_2038;
  assign GEN_2040 = 9'h55 == T_24222 ? T_23676_85 : GEN_2039;
  assign GEN_2041 = 9'h56 == T_24222 ? T_23676_86 : GEN_2040;
  assign GEN_2042 = 9'h57 == T_24222 ? T_23676_87 : GEN_2041;
  assign GEN_2043 = 9'h58 == T_24222 ? T_23676_88 : GEN_2042;
  assign GEN_2044 = 9'h59 == T_24222 ? T_23676_89 : GEN_2043;
  assign GEN_2045 = 9'h5a == T_24222 ? T_23676_90 : GEN_2044;
  assign GEN_2046 = 9'h5b == T_24222 ? T_23676_91 : GEN_2045;
  assign GEN_2047 = 9'h5c == T_24222 ? T_23676_92 : GEN_2046;
  assign GEN_2048 = 9'h5d == T_24222 ? T_23676_93 : GEN_2047;
  assign GEN_2049 = 9'h5e == T_24222 ? T_23676_94 : GEN_2048;
  assign GEN_2050 = 9'h5f == T_24222 ? T_23676_95 : GEN_2049;
  assign GEN_2051 = 9'h60 == T_24222 ? T_23676_96 : GEN_2050;
  assign GEN_2052 = 9'h61 == T_24222 ? T_23676_97 : GEN_2051;
  assign GEN_2053 = 9'h62 == T_24222 ? T_23676_98 : GEN_2052;
  assign GEN_2054 = 9'h63 == T_24222 ? T_23676_99 : GEN_2053;
  assign GEN_2055 = 9'h64 == T_24222 ? T_23676_100 : GEN_2054;
  assign GEN_2056 = 9'h65 == T_24222 ? T_23676_101 : GEN_2055;
  assign GEN_2057 = 9'h66 == T_24222 ? T_23676_102 : GEN_2056;
  assign GEN_2058 = 9'h67 == T_24222 ? T_23676_103 : GEN_2057;
  assign GEN_2059 = 9'h68 == T_24222 ? T_23676_104 : GEN_2058;
  assign GEN_2060 = 9'h69 == T_24222 ? T_23676_105 : GEN_2059;
  assign GEN_2061 = 9'h6a == T_24222 ? T_23676_106 : GEN_2060;
  assign GEN_2062 = 9'h6b == T_24222 ? T_23676_107 : GEN_2061;
  assign GEN_2063 = 9'h6c == T_24222 ? T_23676_108 : GEN_2062;
  assign GEN_2064 = 9'h6d == T_24222 ? T_23676_109 : GEN_2063;
  assign GEN_2065 = 9'h6e == T_24222 ? T_23676_110 : GEN_2064;
  assign GEN_2066 = 9'h6f == T_24222 ? T_23676_111 : GEN_2065;
  assign GEN_2067 = 9'h70 == T_24222 ? T_23676_112 : GEN_2066;
  assign GEN_2068 = 9'h71 == T_24222 ? T_23676_113 : GEN_2067;
  assign GEN_2069 = 9'h72 == T_24222 ? T_23676_114 : GEN_2068;
  assign GEN_2070 = 9'h73 == T_24222 ? T_23676_115 : GEN_2069;
  assign GEN_2071 = 9'h74 == T_24222 ? T_23676_116 : GEN_2070;
  assign GEN_2072 = 9'h75 == T_24222 ? T_23676_117 : GEN_2071;
  assign GEN_2073 = 9'h76 == T_24222 ? T_23676_118 : GEN_2072;
  assign GEN_2074 = 9'h77 == T_24222 ? T_23676_119 : GEN_2073;
  assign GEN_2075 = 9'h78 == T_24222 ? T_23676_120 : GEN_2074;
  assign GEN_2076 = 9'h79 == T_24222 ? T_23676_121 : GEN_2075;
  assign GEN_2077 = 9'h7a == T_24222 ? T_23676_122 : GEN_2076;
  assign GEN_2078 = 9'h7b == T_24222 ? T_23676_123 : GEN_2077;
  assign GEN_2079 = 9'h7c == T_24222 ? T_23676_124 : GEN_2078;
  assign GEN_2080 = 9'h7d == T_24222 ? T_23676_125 : GEN_2079;
  assign GEN_2081 = 9'h7e == T_24222 ? T_23676_126 : GEN_2080;
  assign GEN_2082 = 9'h7f == T_24222 ? T_23676_127 : GEN_2081;
  assign GEN_2083 = 9'h80 == T_24222 ? T_23676_128 : GEN_2082;
  assign GEN_2084 = 9'h81 == T_24222 ? T_23676_129 : GEN_2083;
  assign GEN_2085 = 9'h82 == T_24222 ? T_23676_130 : GEN_2084;
  assign GEN_2086 = 9'h83 == T_24222 ? T_23676_131 : GEN_2085;
  assign GEN_2087 = 9'h84 == T_24222 ? T_23676_132 : GEN_2086;
  assign GEN_2088 = 9'h85 == T_24222 ? T_23676_133 : GEN_2087;
  assign GEN_2089 = 9'h86 == T_24222 ? T_23676_134 : GEN_2088;
  assign GEN_2090 = 9'h87 == T_24222 ? T_23676_135 : GEN_2089;
  assign GEN_2091 = 9'h88 == T_24222 ? T_23676_136 : GEN_2090;
  assign GEN_2092 = 9'h89 == T_24222 ? T_23676_137 : GEN_2091;
  assign GEN_2093 = 9'h8a == T_24222 ? T_23676_138 : GEN_2092;
  assign GEN_2094 = 9'h8b == T_24222 ? T_23676_139 : GEN_2093;
  assign GEN_2095 = 9'h8c == T_24222 ? T_23676_140 : GEN_2094;
  assign GEN_2096 = 9'h8d == T_24222 ? T_23676_141 : GEN_2095;
  assign GEN_2097 = 9'h8e == T_24222 ? T_23676_142 : GEN_2096;
  assign GEN_2098 = 9'h8f == T_24222 ? T_23676_143 : GEN_2097;
  assign GEN_2099 = 9'h90 == T_24222 ? T_23676_144 : GEN_2098;
  assign GEN_2100 = 9'h91 == T_24222 ? T_23676_145 : GEN_2099;
  assign GEN_2101 = 9'h92 == T_24222 ? T_23676_146 : GEN_2100;
  assign GEN_2102 = 9'h93 == T_24222 ? T_23676_147 : GEN_2101;
  assign GEN_2103 = 9'h94 == T_24222 ? T_23676_148 : GEN_2102;
  assign GEN_2104 = 9'h95 == T_24222 ? T_23676_149 : GEN_2103;
  assign GEN_2105 = 9'h96 == T_24222 ? T_23676_150 : GEN_2104;
  assign GEN_2106 = 9'h97 == T_24222 ? T_23676_151 : GEN_2105;
  assign GEN_2107 = 9'h98 == T_24222 ? T_23676_152 : GEN_2106;
  assign GEN_2108 = 9'h99 == T_24222 ? T_23676_153 : GEN_2107;
  assign GEN_2109 = 9'h9a == T_24222 ? T_23676_154 : GEN_2108;
  assign GEN_2110 = 9'h9b == T_24222 ? T_23676_155 : GEN_2109;
  assign GEN_2111 = 9'h9c == T_24222 ? T_23676_156 : GEN_2110;
  assign GEN_2112 = 9'h9d == T_24222 ? T_23676_157 : GEN_2111;
  assign GEN_2113 = 9'h9e == T_24222 ? T_23676_158 : GEN_2112;
  assign GEN_2114 = 9'h9f == T_24222 ? T_23676_159 : GEN_2113;
  assign GEN_2115 = 9'ha0 == T_24222 ? T_23676_160 : GEN_2114;
  assign GEN_2116 = 9'ha1 == T_24222 ? T_23676_161 : GEN_2115;
  assign GEN_2117 = 9'ha2 == T_24222 ? T_23676_162 : GEN_2116;
  assign GEN_2118 = 9'ha3 == T_24222 ? T_23676_163 : GEN_2117;
  assign GEN_2119 = 9'ha4 == T_24222 ? T_23676_164 : GEN_2118;
  assign GEN_2120 = 9'ha5 == T_24222 ? T_23676_165 : GEN_2119;
  assign GEN_2121 = 9'ha6 == T_24222 ? T_23676_166 : GEN_2120;
  assign GEN_2122 = 9'ha7 == T_24222 ? T_23676_167 : GEN_2121;
  assign GEN_2123 = 9'ha8 == T_24222 ? T_23676_168 : GEN_2122;
  assign GEN_2124 = 9'ha9 == T_24222 ? T_23676_169 : GEN_2123;
  assign GEN_2125 = 9'haa == T_24222 ? T_23676_170 : GEN_2124;
  assign GEN_2126 = 9'hab == T_24222 ? T_23676_171 : GEN_2125;
  assign GEN_2127 = 9'hac == T_24222 ? T_23676_172 : GEN_2126;
  assign GEN_2128 = 9'had == T_24222 ? T_23676_173 : GEN_2127;
  assign GEN_2129 = 9'hae == T_24222 ? T_23676_174 : GEN_2128;
  assign GEN_2130 = 9'haf == T_24222 ? T_23676_175 : GEN_2129;
  assign GEN_2131 = 9'hb0 == T_24222 ? T_23676_176 : GEN_2130;
  assign GEN_2132 = 9'hb1 == T_24222 ? T_23676_177 : GEN_2131;
  assign GEN_2133 = 9'hb2 == T_24222 ? T_23676_178 : GEN_2132;
  assign GEN_2134 = 9'hb3 == T_24222 ? T_23676_179 : GEN_2133;
  assign GEN_2135 = 9'hb4 == T_24222 ? T_23676_180 : GEN_2134;
  assign GEN_2136 = 9'hb5 == T_24222 ? T_23676_181 : GEN_2135;
  assign GEN_2137 = 9'hb6 == T_24222 ? T_23676_182 : GEN_2136;
  assign GEN_2138 = 9'hb7 == T_24222 ? T_23676_183 : GEN_2137;
  assign GEN_2139 = 9'hb8 == T_24222 ? T_23676_184 : GEN_2138;
  assign GEN_2140 = 9'hb9 == T_24222 ? T_23676_185 : GEN_2139;
  assign GEN_2141 = 9'hba == T_24222 ? T_23676_186 : GEN_2140;
  assign GEN_2142 = 9'hbb == T_24222 ? T_23676_187 : GEN_2141;
  assign GEN_2143 = 9'hbc == T_24222 ? T_23676_188 : GEN_2142;
  assign GEN_2144 = 9'hbd == T_24222 ? T_23676_189 : GEN_2143;
  assign GEN_2145 = 9'hbe == T_24222 ? T_23676_190 : GEN_2144;
  assign GEN_2146 = 9'hbf == T_24222 ? T_23676_191 : GEN_2145;
  assign GEN_2147 = 9'hc0 == T_24222 ? T_23676_192 : GEN_2146;
  assign GEN_2148 = 9'hc1 == T_24222 ? T_23676_193 : GEN_2147;
  assign GEN_2149 = 9'hc2 == T_24222 ? T_23676_194 : GEN_2148;
  assign GEN_2150 = 9'hc3 == T_24222 ? T_23676_195 : GEN_2149;
  assign GEN_2151 = 9'hc4 == T_24222 ? T_23676_196 : GEN_2150;
  assign GEN_2152 = 9'hc5 == T_24222 ? T_23676_197 : GEN_2151;
  assign GEN_2153 = 9'hc6 == T_24222 ? T_23676_198 : GEN_2152;
  assign GEN_2154 = 9'hc7 == T_24222 ? T_23676_199 : GEN_2153;
  assign GEN_2155 = 9'hc8 == T_24222 ? T_23676_200 : GEN_2154;
  assign GEN_2156 = 9'hc9 == T_24222 ? T_23676_201 : GEN_2155;
  assign GEN_2157 = 9'hca == T_24222 ? T_23676_202 : GEN_2156;
  assign GEN_2158 = 9'hcb == T_24222 ? T_23676_203 : GEN_2157;
  assign GEN_2159 = 9'hcc == T_24222 ? T_23676_204 : GEN_2158;
  assign GEN_2160 = 9'hcd == T_24222 ? T_23676_205 : GEN_2159;
  assign GEN_2161 = 9'hce == T_24222 ? T_23676_206 : GEN_2160;
  assign GEN_2162 = 9'hcf == T_24222 ? T_23676_207 : GEN_2161;
  assign GEN_2163 = 9'hd0 == T_24222 ? T_23676_208 : GEN_2162;
  assign GEN_2164 = 9'hd1 == T_24222 ? T_23676_209 : GEN_2163;
  assign GEN_2165 = 9'hd2 == T_24222 ? T_23676_210 : GEN_2164;
  assign GEN_2166 = 9'hd3 == T_24222 ? T_23676_211 : GEN_2165;
  assign GEN_2167 = 9'hd4 == T_24222 ? T_23676_212 : GEN_2166;
  assign GEN_2168 = 9'hd5 == T_24222 ? T_23676_213 : GEN_2167;
  assign GEN_2169 = 9'hd6 == T_24222 ? T_23676_214 : GEN_2168;
  assign GEN_2170 = 9'hd7 == T_24222 ? T_23676_215 : GEN_2169;
  assign GEN_2171 = 9'hd8 == T_24222 ? T_23676_216 : GEN_2170;
  assign GEN_2172 = 9'hd9 == T_24222 ? T_23676_217 : GEN_2171;
  assign GEN_2173 = 9'hda == T_24222 ? T_23676_218 : GEN_2172;
  assign GEN_2174 = 9'hdb == T_24222 ? T_23676_219 : GEN_2173;
  assign GEN_2175 = 9'hdc == T_24222 ? T_23676_220 : GEN_2174;
  assign GEN_2176 = 9'hdd == T_24222 ? T_23676_221 : GEN_2175;
  assign GEN_2177 = 9'hde == T_24222 ? T_23676_222 : GEN_2176;
  assign GEN_2178 = 9'hdf == T_24222 ? T_23676_223 : GEN_2177;
  assign GEN_2179 = 9'he0 == T_24222 ? T_23676_224 : GEN_2178;
  assign GEN_2180 = 9'he1 == T_24222 ? T_23676_225 : GEN_2179;
  assign GEN_2181 = 9'he2 == T_24222 ? T_23676_226 : GEN_2180;
  assign GEN_2182 = 9'he3 == T_24222 ? T_23676_227 : GEN_2181;
  assign GEN_2183 = 9'he4 == T_24222 ? T_23676_228 : GEN_2182;
  assign GEN_2184 = 9'he5 == T_24222 ? T_23676_229 : GEN_2183;
  assign GEN_2185 = 9'he6 == T_24222 ? T_23676_230 : GEN_2184;
  assign GEN_2186 = 9'he7 == T_24222 ? T_23676_231 : GEN_2185;
  assign GEN_2187 = 9'he8 == T_24222 ? T_23676_232 : GEN_2186;
  assign GEN_2188 = 9'he9 == T_24222 ? T_23676_233 : GEN_2187;
  assign GEN_2189 = 9'hea == T_24222 ? T_23676_234 : GEN_2188;
  assign GEN_2190 = 9'heb == T_24222 ? T_23676_235 : GEN_2189;
  assign GEN_2191 = 9'hec == T_24222 ? T_23676_236 : GEN_2190;
  assign GEN_2192 = 9'hed == T_24222 ? T_23676_237 : GEN_2191;
  assign GEN_2193 = 9'hee == T_24222 ? T_23676_238 : GEN_2192;
  assign GEN_2194 = 9'hef == T_24222 ? T_23676_239 : GEN_2193;
  assign GEN_2195 = 9'hf0 == T_24222 ? T_23676_240 : GEN_2194;
  assign GEN_2196 = 9'hf1 == T_24222 ? T_23676_241 : GEN_2195;
  assign GEN_2197 = 9'hf2 == T_24222 ? T_23676_242 : GEN_2196;
  assign GEN_2198 = 9'hf3 == T_24222 ? T_23676_243 : GEN_2197;
  assign GEN_2199 = 9'hf4 == T_24222 ? T_23676_244 : GEN_2198;
  assign GEN_2200 = 9'hf5 == T_24222 ? T_23676_245 : GEN_2199;
  assign GEN_2201 = 9'hf6 == T_24222 ? T_23676_246 : GEN_2200;
  assign GEN_2202 = 9'hf7 == T_24222 ? T_23676_247 : GEN_2201;
  assign GEN_2203 = 9'hf8 == T_24222 ? T_23676_248 : GEN_2202;
  assign GEN_2204 = 9'hf9 == T_24222 ? T_23676_249 : GEN_2203;
  assign GEN_2205 = 9'hfa == T_24222 ? T_23676_250 : GEN_2204;
  assign GEN_2206 = 9'hfb == T_24222 ? T_23676_251 : GEN_2205;
  assign GEN_2207 = 9'hfc == T_24222 ? T_23676_252 : GEN_2206;
  assign GEN_2208 = 9'hfd == T_24222 ? T_23676_253 : GEN_2207;
  assign GEN_2209 = 9'hfe == T_24222 ? T_23676_254 : GEN_2208;
  assign GEN_2210 = 9'hff == T_24222 ? T_23676_255 : GEN_2209;
  assign GEN_2211 = 9'h100 == T_24222 ? T_23676_256 : GEN_2210;
  assign GEN_2212 = 9'h101 == T_24222 ? T_23676_257 : GEN_2211;
  assign GEN_2213 = 9'h102 == T_24222 ? T_23676_258 : GEN_2212;
  assign GEN_2214 = 9'h103 == T_24222 ? T_23676_259 : GEN_2213;
  assign GEN_2215 = 9'h104 == T_24222 ? T_23676_260 : GEN_2214;
  assign GEN_2216 = 9'h105 == T_24222 ? T_23676_261 : GEN_2215;
  assign GEN_2217 = 9'h106 == T_24222 ? T_23676_262 : GEN_2216;
  assign GEN_2218 = 9'h107 == T_24222 ? T_23676_263 : GEN_2217;
  assign GEN_2219 = 9'h108 == T_24222 ? T_23676_264 : GEN_2218;
  assign GEN_2220 = 9'h109 == T_24222 ? T_23676_265 : GEN_2219;
  assign GEN_2221 = 9'h10a == T_24222 ? T_23676_266 : GEN_2220;
  assign GEN_2222 = 9'h10b == T_24222 ? T_23676_267 : GEN_2221;
  assign GEN_2223 = 9'h10c == T_24222 ? T_23676_268 : GEN_2222;
  assign GEN_2224 = 9'h10d == T_24222 ? T_23676_269 : GEN_2223;
  assign GEN_2225 = 9'h10e == T_24222 ? T_23676_270 : GEN_2224;
  assign GEN_2226 = 9'h10f == T_24222 ? T_23676_271 : GEN_2225;
  assign GEN_2227 = 9'h110 == T_24222 ? T_23676_272 : GEN_2226;
  assign GEN_2228 = 9'h111 == T_24222 ? T_23676_273 : GEN_2227;
  assign GEN_2229 = 9'h112 == T_24222 ? T_23676_274 : GEN_2228;
  assign GEN_2230 = 9'h113 == T_24222 ? T_23676_275 : GEN_2229;
  assign GEN_2231 = 9'h114 == T_24222 ? T_23676_276 : GEN_2230;
  assign GEN_2232 = 9'h115 == T_24222 ? T_23676_277 : GEN_2231;
  assign GEN_2233 = 9'h116 == T_24222 ? T_23676_278 : GEN_2232;
  assign GEN_2234 = 9'h117 == T_24222 ? T_23676_279 : GEN_2233;
  assign GEN_2235 = 9'h118 == T_24222 ? T_23676_280 : GEN_2234;
  assign GEN_2236 = 9'h119 == T_24222 ? T_23676_281 : GEN_2235;
  assign GEN_2237 = 9'h11a == T_24222 ? T_23676_282 : GEN_2236;
  assign GEN_2238 = 9'h11b == T_24222 ? T_23676_283 : GEN_2237;
  assign GEN_2239 = 9'h11c == T_24222 ? T_23676_284 : GEN_2238;
  assign GEN_2240 = 9'h11d == T_24222 ? T_23676_285 : GEN_2239;
  assign GEN_2241 = 9'h11e == T_24222 ? T_23676_286 : GEN_2240;
  assign GEN_2242 = 9'h11f == T_24222 ? T_23676_287 : GEN_2241;
  assign GEN_2243 = 9'h120 == T_24222 ? T_23676_288 : GEN_2242;
  assign GEN_2244 = 9'h121 == T_24222 ? T_23676_289 : GEN_2243;
  assign GEN_2245 = 9'h122 == T_24222 ? T_23676_290 : GEN_2244;
  assign GEN_2246 = 9'h123 == T_24222 ? T_23676_291 : GEN_2245;
  assign GEN_2247 = 9'h124 == T_24222 ? T_23676_292 : GEN_2246;
  assign GEN_2248 = 9'h125 == T_24222 ? T_23676_293 : GEN_2247;
  assign GEN_2249 = 9'h126 == T_24222 ? T_23676_294 : GEN_2248;
  assign GEN_2250 = 9'h127 == T_24222 ? T_23676_295 : GEN_2249;
  assign GEN_2251 = 9'h128 == T_24222 ? T_23676_296 : GEN_2250;
  assign GEN_2252 = 9'h129 == T_24222 ? T_23676_297 : GEN_2251;
  assign GEN_2253 = 9'h12a == T_24222 ? T_23676_298 : GEN_2252;
  assign GEN_2254 = 9'h12b == T_24222 ? T_23676_299 : GEN_2253;
  assign GEN_2255 = 9'h12c == T_24222 ? T_23676_300 : GEN_2254;
  assign GEN_2256 = 9'h12d == T_24222 ? T_23676_301 : GEN_2255;
  assign GEN_2257 = 9'h12e == T_24222 ? T_23676_302 : GEN_2256;
  assign GEN_2258 = 9'h12f == T_24222 ? T_23676_303 : GEN_2257;
  assign GEN_2259 = 9'h130 == T_24222 ? T_23676_304 : GEN_2258;
  assign GEN_2260 = 9'h131 == T_24222 ? T_23676_305 : GEN_2259;
  assign GEN_2261 = 9'h132 == T_24222 ? T_23676_306 : GEN_2260;
  assign GEN_2262 = 9'h133 == T_24222 ? T_23676_307 : GEN_2261;
  assign GEN_2263 = 9'h134 == T_24222 ? T_23676_308 : GEN_2262;
  assign GEN_2264 = 9'h135 == T_24222 ? T_23676_309 : GEN_2263;
  assign GEN_2265 = 9'h136 == T_24222 ? T_23676_310 : GEN_2264;
  assign GEN_2266 = 9'h137 == T_24222 ? T_23676_311 : GEN_2265;
  assign GEN_2267 = 9'h138 == T_24222 ? T_23676_312 : GEN_2266;
  assign GEN_2268 = 9'h139 == T_24222 ? T_23676_313 : GEN_2267;
  assign GEN_2269 = 9'h13a == T_24222 ? T_23676_314 : GEN_2268;
  assign GEN_2270 = 9'h13b == T_24222 ? T_23676_315 : GEN_2269;
  assign GEN_2271 = 9'h13c == T_24222 ? T_23676_316 : GEN_2270;
  assign GEN_2272 = 9'h13d == T_24222 ? T_23676_317 : GEN_2271;
  assign GEN_2273 = 9'h13e == T_24222 ? T_23676_318 : GEN_2272;
  assign GEN_2274 = 9'h13f == T_24222 ? T_23676_319 : GEN_2273;
  assign GEN_2275 = 9'h140 == T_24222 ? T_23676_320 : GEN_2274;
  assign GEN_2276 = 9'h141 == T_24222 ? T_23676_321 : GEN_2275;
  assign GEN_2277 = 9'h142 == T_24222 ? T_23676_322 : GEN_2276;
  assign GEN_2278 = 9'h143 == T_24222 ? T_23676_323 : GEN_2277;
  assign GEN_2279 = 9'h144 == T_24222 ? T_23676_324 : GEN_2278;
  assign GEN_2280 = 9'h145 == T_24222 ? T_23676_325 : GEN_2279;
  assign GEN_2281 = 9'h146 == T_24222 ? T_23676_326 : GEN_2280;
  assign GEN_2282 = 9'h147 == T_24222 ? T_23676_327 : GEN_2281;
  assign GEN_2283 = 9'h148 == T_24222 ? T_23676_328 : GEN_2282;
  assign GEN_2284 = 9'h149 == T_24222 ? T_23676_329 : GEN_2283;
  assign GEN_2285 = 9'h14a == T_24222 ? T_23676_330 : GEN_2284;
  assign GEN_2286 = 9'h14b == T_24222 ? T_23676_331 : GEN_2285;
  assign GEN_2287 = 9'h14c == T_24222 ? T_23676_332 : GEN_2286;
  assign GEN_2288 = 9'h14d == T_24222 ? T_23676_333 : GEN_2287;
  assign GEN_2289 = 9'h14e == T_24222 ? T_23676_334 : GEN_2288;
  assign GEN_2290 = 9'h14f == T_24222 ? T_23676_335 : GEN_2289;
  assign GEN_2291 = 9'h150 == T_24222 ? T_23676_336 : GEN_2290;
  assign GEN_2292 = 9'h151 == T_24222 ? T_23676_337 : GEN_2291;
  assign GEN_2293 = 9'h152 == T_24222 ? T_23676_338 : GEN_2292;
  assign GEN_2294 = 9'h153 == T_24222 ? T_23676_339 : GEN_2293;
  assign GEN_2295 = 9'h154 == T_24222 ? T_23676_340 : GEN_2294;
  assign GEN_2296 = 9'h155 == T_24222 ? T_23676_341 : GEN_2295;
  assign GEN_2297 = 9'h156 == T_24222 ? T_23676_342 : GEN_2296;
  assign GEN_2298 = 9'h157 == T_24222 ? T_23676_343 : GEN_2297;
  assign GEN_2299 = 9'h158 == T_24222 ? T_23676_344 : GEN_2298;
  assign GEN_2300 = 9'h159 == T_24222 ? T_23676_345 : GEN_2299;
  assign GEN_2301 = 9'h15a == T_24222 ? T_23676_346 : GEN_2300;
  assign GEN_2302 = 9'h15b == T_24222 ? T_23676_347 : GEN_2301;
  assign GEN_2303 = 9'h15c == T_24222 ? T_23676_348 : GEN_2302;
  assign GEN_2304 = 9'h15d == T_24222 ? T_23676_349 : GEN_2303;
  assign GEN_2305 = 9'h15e == T_24222 ? T_23676_350 : GEN_2304;
  assign GEN_2306 = 9'h15f == T_24222 ? T_23676_351 : GEN_2305;
  assign GEN_2307 = 9'h160 == T_24222 ? T_23676_352 : GEN_2306;
  assign GEN_2308 = 9'h161 == T_24222 ? T_23676_353 : GEN_2307;
  assign GEN_2309 = 9'h162 == T_24222 ? T_23676_354 : GEN_2308;
  assign GEN_2310 = 9'h163 == T_24222 ? T_23676_355 : GEN_2309;
  assign GEN_2311 = 9'h164 == T_24222 ? T_23676_356 : GEN_2310;
  assign GEN_2312 = 9'h165 == T_24222 ? T_23676_357 : GEN_2311;
  assign GEN_2313 = 9'h166 == T_24222 ? T_23676_358 : GEN_2312;
  assign GEN_2314 = 9'h167 == T_24222 ? T_23676_359 : GEN_2313;
  assign GEN_2315 = 9'h168 == T_24222 ? T_23676_360 : GEN_2314;
  assign GEN_2316 = 9'h169 == T_24222 ? T_23676_361 : GEN_2315;
  assign GEN_2317 = 9'h16a == T_24222 ? T_23676_362 : GEN_2316;
  assign GEN_2318 = 9'h16b == T_24222 ? T_23676_363 : GEN_2317;
  assign GEN_2319 = 9'h16c == T_24222 ? T_23676_364 : GEN_2318;
  assign GEN_2320 = 9'h16d == T_24222 ? T_23676_365 : GEN_2319;
  assign GEN_2321 = 9'h16e == T_24222 ? T_23676_366 : GEN_2320;
  assign GEN_2322 = 9'h16f == T_24222 ? T_23676_367 : GEN_2321;
  assign GEN_2323 = 9'h170 == T_24222 ? T_23676_368 : GEN_2322;
  assign GEN_2324 = 9'h171 == T_24222 ? T_23676_369 : GEN_2323;
  assign GEN_2325 = 9'h172 == T_24222 ? T_23676_370 : GEN_2324;
  assign GEN_2326 = 9'h173 == T_24222 ? T_23676_371 : GEN_2325;
  assign GEN_2327 = 9'h174 == T_24222 ? T_23676_372 : GEN_2326;
  assign GEN_2328 = 9'h175 == T_24222 ? T_23676_373 : GEN_2327;
  assign GEN_2329 = 9'h176 == T_24222 ? T_23676_374 : GEN_2328;
  assign GEN_2330 = 9'h177 == T_24222 ? T_23676_375 : GEN_2329;
  assign GEN_2331 = 9'h178 == T_24222 ? T_23676_376 : GEN_2330;
  assign GEN_2332 = 9'h179 == T_24222 ? T_23676_377 : GEN_2331;
  assign GEN_2333 = 9'h17a == T_24222 ? T_23676_378 : GEN_2332;
  assign GEN_2334 = 9'h17b == T_24222 ? T_23676_379 : GEN_2333;
  assign GEN_2335 = 9'h17c == T_24222 ? T_23676_380 : GEN_2334;
  assign GEN_2336 = 9'h17d == T_24222 ? T_23676_381 : GEN_2335;
  assign GEN_2337 = 9'h17e == T_24222 ? T_23676_382 : GEN_2336;
  assign GEN_2338 = 9'h17f == T_24222 ? T_23676_383 : GEN_2337;
  assign GEN_2339 = 9'h180 == T_24222 ? T_23676_384 : GEN_2338;
  assign GEN_2340 = 9'h181 == T_24222 ? T_23676_385 : GEN_2339;
  assign GEN_2341 = 9'h182 == T_24222 ? T_23676_386 : GEN_2340;
  assign GEN_2342 = 9'h183 == T_24222 ? T_23676_387 : GEN_2341;
  assign GEN_2343 = 9'h184 == T_24222 ? T_23676_388 : GEN_2342;
  assign GEN_2344 = 9'h185 == T_24222 ? T_23676_389 : GEN_2343;
  assign GEN_2345 = 9'h186 == T_24222 ? T_23676_390 : GEN_2344;
  assign GEN_2346 = 9'h187 == T_24222 ? T_23676_391 : GEN_2345;
  assign GEN_2347 = 9'h188 == T_24222 ? T_23676_392 : GEN_2346;
  assign GEN_2348 = 9'h189 == T_24222 ? T_23676_393 : GEN_2347;
  assign GEN_2349 = 9'h18a == T_24222 ? T_23676_394 : GEN_2348;
  assign GEN_2350 = 9'h18b == T_24222 ? T_23676_395 : GEN_2349;
  assign GEN_2351 = 9'h18c == T_24222 ? T_23676_396 : GEN_2350;
  assign GEN_2352 = 9'h18d == T_24222 ? T_23676_397 : GEN_2351;
  assign GEN_2353 = 9'h18e == T_24222 ? T_23676_398 : GEN_2352;
  assign GEN_2354 = 9'h18f == T_24222 ? T_23676_399 : GEN_2353;
  assign GEN_2355 = 9'h190 == T_24222 ? T_23676_400 : GEN_2354;
  assign GEN_2356 = 9'h191 == T_24222 ? T_23676_401 : GEN_2355;
  assign GEN_2357 = 9'h192 == T_24222 ? T_23676_402 : GEN_2356;
  assign GEN_2358 = 9'h193 == T_24222 ? T_23676_403 : GEN_2357;
  assign GEN_2359 = 9'h194 == T_24222 ? T_23676_404 : GEN_2358;
  assign GEN_2360 = 9'h195 == T_24222 ? T_23676_405 : GEN_2359;
  assign GEN_2361 = 9'h196 == T_24222 ? T_23676_406 : GEN_2360;
  assign GEN_2362 = 9'h197 == T_24222 ? T_23676_407 : GEN_2361;
  assign GEN_2363 = 9'h198 == T_24222 ? T_23676_408 : GEN_2362;
  assign GEN_2364 = 9'h199 == T_24222 ? T_23676_409 : GEN_2363;
  assign GEN_2365 = 9'h19a == T_24222 ? T_23676_410 : GEN_2364;
  assign GEN_2366 = 9'h19b == T_24222 ? T_23676_411 : GEN_2365;
  assign GEN_2367 = 9'h19c == T_24222 ? T_23676_412 : GEN_2366;
  assign GEN_2368 = 9'h19d == T_24222 ? T_23676_413 : GEN_2367;
  assign GEN_2369 = 9'h19e == T_24222 ? T_23676_414 : GEN_2368;
  assign GEN_2370 = 9'h19f == T_24222 ? T_23676_415 : GEN_2369;
  assign GEN_2371 = 9'h1a0 == T_24222 ? T_23676_416 : GEN_2370;
  assign GEN_2372 = 9'h1a1 == T_24222 ? T_23676_417 : GEN_2371;
  assign GEN_2373 = 9'h1a2 == T_24222 ? T_23676_418 : GEN_2372;
  assign GEN_2374 = 9'h1a3 == T_24222 ? T_23676_419 : GEN_2373;
  assign GEN_2375 = 9'h1a4 == T_24222 ? T_23676_420 : GEN_2374;
  assign GEN_2376 = 9'h1a5 == T_24222 ? T_23676_421 : GEN_2375;
  assign GEN_2377 = 9'h1a6 == T_24222 ? T_23676_422 : GEN_2376;
  assign GEN_2378 = 9'h1a7 == T_24222 ? T_23676_423 : GEN_2377;
  assign GEN_2379 = 9'h1a8 == T_24222 ? T_23676_424 : GEN_2378;
  assign GEN_2380 = 9'h1a9 == T_24222 ? T_23676_425 : GEN_2379;
  assign GEN_2381 = 9'h1aa == T_24222 ? T_23676_426 : GEN_2380;
  assign GEN_2382 = 9'h1ab == T_24222 ? T_23676_427 : GEN_2381;
  assign GEN_2383 = 9'h1ac == T_24222 ? T_23676_428 : GEN_2382;
  assign GEN_2384 = 9'h1ad == T_24222 ? T_23676_429 : GEN_2383;
  assign GEN_2385 = 9'h1ae == T_24222 ? T_23676_430 : GEN_2384;
  assign GEN_2386 = 9'h1af == T_24222 ? T_23676_431 : GEN_2385;
  assign GEN_2387 = 9'h1b0 == T_24222 ? T_23676_432 : GEN_2386;
  assign GEN_2388 = 9'h1b1 == T_24222 ? T_23676_433 : GEN_2387;
  assign GEN_2389 = 9'h1b2 == T_24222 ? T_23676_434 : GEN_2388;
  assign GEN_2390 = 9'h1b3 == T_24222 ? T_23676_435 : GEN_2389;
  assign GEN_2391 = 9'h1b4 == T_24222 ? T_23676_436 : GEN_2390;
  assign GEN_2392 = 9'h1b5 == T_24222 ? T_23676_437 : GEN_2391;
  assign GEN_2393 = 9'h1b6 == T_24222 ? T_23676_438 : GEN_2392;
  assign GEN_2394 = 9'h1b7 == T_24222 ? T_23676_439 : GEN_2393;
  assign GEN_2395 = 9'h1b8 == T_24222 ? T_23676_440 : GEN_2394;
  assign GEN_2396 = 9'h1b9 == T_24222 ? T_23676_441 : GEN_2395;
  assign GEN_2397 = 9'h1ba == T_24222 ? T_23676_442 : GEN_2396;
  assign GEN_2398 = 9'h1bb == T_24222 ? T_23676_443 : GEN_2397;
  assign GEN_2399 = 9'h1bc == T_24222 ? T_23676_444 : GEN_2398;
  assign GEN_2400 = 9'h1bd == T_24222 ? T_23676_445 : GEN_2399;
  assign GEN_2401 = 9'h1be == T_24222 ? T_23676_446 : GEN_2400;
  assign GEN_2402 = 9'h1bf == T_24222 ? T_23676_447 : GEN_2401;
  assign GEN_2403 = 9'h1c0 == T_24222 ? T_23676_448 : GEN_2402;
  assign GEN_2404 = 9'h1c1 == T_24222 ? T_23676_449 : GEN_2403;
  assign GEN_2405 = 9'h1c2 == T_24222 ? T_23676_450 : GEN_2404;
  assign GEN_2406 = 9'h1c3 == T_24222 ? T_23676_451 : GEN_2405;
  assign GEN_2407 = 9'h1c4 == T_24222 ? T_23676_452 : GEN_2406;
  assign GEN_2408 = 9'h1c5 == T_24222 ? T_23676_453 : GEN_2407;
  assign GEN_2409 = 9'h1c6 == T_24222 ? T_23676_454 : GEN_2408;
  assign GEN_2410 = 9'h1c7 == T_24222 ? T_23676_455 : GEN_2409;
  assign GEN_2411 = 9'h1c8 == T_24222 ? T_23676_456 : GEN_2410;
  assign GEN_2412 = 9'h1c9 == T_24222 ? T_23676_457 : GEN_2411;
  assign GEN_2413 = 9'h1ca == T_24222 ? T_23676_458 : GEN_2412;
  assign GEN_2414 = 9'h1cb == T_24222 ? T_23676_459 : GEN_2413;
  assign GEN_2415 = 9'h1cc == T_24222 ? T_23676_460 : GEN_2414;
  assign GEN_2416 = 9'h1cd == T_24222 ? T_23676_461 : GEN_2415;
  assign GEN_2417 = 9'h1ce == T_24222 ? T_23676_462 : GEN_2416;
  assign GEN_2418 = 9'h1cf == T_24222 ? T_23676_463 : GEN_2417;
  assign GEN_2419 = 9'h1d0 == T_24222 ? T_23676_464 : GEN_2418;
  assign GEN_2420 = 9'h1d1 == T_24222 ? T_23676_465 : GEN_2419;
  assign GEN_2421 = 9'h1d2 == T_24222 ? T_23676_466 : GEN_2420;
  assign GEN_2422 = 9'h1d3 == T_24222 ? T_23676_467 : GEN_2421;
  assign GEN_2423 = 9'h1d4 == T_24222 ? T_23676_468 : GEN_2422;
  assign GEN_2424 = 9'h1d5 == T_24222 ? T_23676_469 : GEN_2423;
  assign GEN_2425 = 9'h1d6 == T_24222 ? T_23676_470 : GEN_2424;
  assign GEN_2426 = 9'h1d7 == T_24222 ? T_23676_471 : GEN_2425;
  assign GEN_2427 = 9'h1d8 == T_24222 ? T_23676_472 : GEN_2426;
  assign GEN_2428 = 9'h1d9 == T_24222 ? T_23676_473 : GEN_2427;
  assign GEN_2429 = 9'h1da == T_24222 ? T_23676_474 : GEN_2428;
  assign GEN_2430 = 9'h1db == T_24222 ? T_23676_475 : GEN_2429;
  assign GEN_2431 = 9'h1dc == T_24222 ? T_23676_476 : GEN_2430;
  assign GEN_2432 = 9'h1dd == T_24222 ? T_23676_477 : GEN_2431;
  assign GEN_2433 = 9'h1de == T_24222 ? T_23676_478 : GEN_2432;
  assign GEN_2434 = 9'h1df == T_24222 ? T_23676_479 : GEN_2433;
  assign GEN_2435 = 9'h1e0 == T_24222 ? T_23676_480 : GEN_2434;
  assign GEN_2436 = 9'h1e1 == T_24222 ? T_23676_481 : GEN_2435;
  assign GEN_2437 = 9'h1e2 == T_24222 ? T_23676_482 : GEN_2436;
  assign GEN_2438 = 9'h1e3 == T_24222 ? T_23676_483 : GEN_2437;
  assign GEN_2439 = 9'h1e4 == T_24222 ? T_23676_484 : GEN_2438;
  assign GEN_2440 = 9'h1e5 == T_24222 ? T_23676_485 : GEN_2439;
  assign GEN_2441 = 9'h1e6 == T_24222 ? T_23676_486 : GEN_2440;
  assign GEN_2442 = 9'h1e7 == T_24222 ? T_23676_487 : GEN_2441;
  assign GEN_2443 = 9'h1e8 == T_24222 ? T_23676_488 : GEN_2442;
  assign GEN_2444 = 9'h1e9 == T_24222 ? T_23676_489 : GEN_2443;
  assign GEN_2445 = 9'h1ea == T_24222 ? T_23676_490 : GEN_2444;
  assign GEN_2446 = 9'h1eb == T_24222 ? T_23676_491 : GEN_2445;
  assign GEN_2447 = 9'h1ec == T_24222 ? T_23676_492 : GEN_2446;
  assign GEN_2448 = 9'h1ed == T_24222 ? T_23676_493 : GEN_2447;
  assign GEN_2449 = 9'h1ee == T_24222 ? T_23676_494 : GEN_2448;
  assign GEN_2450 = 9'h1ef == T_24222 ? T_23676_495 : GEN_2449;
  assign GEN_2451 = 9'h1f0 == T_24222 ? T_23676_496 : GEN_2450;
  assign GEN_2452 = 9'h1f1 == T_24222 ? T_23676_497 : GEN_2451;
  assign GEN_2453 = 9'h1f2 == T_24222 ? T_23676_498 : GEN_2452;
  assign GEN_2454 = 9'h1f3 == T_24222 ? T_23676_499 : GEN_2453;
  assign GEN_2455 = 9'h1f4 == T_24222 ? T_23676_500 : GEN_2454;
  assign GEN_2456 = 9'h1f5 == T_24222 ? T_23676_501 : GEN_2455;
  assign GEN_2457 = 9'h1f6 == T_24222 ? T_23676_502 : GEN_2456;
  assign GEN_2458 = 9'h1f7 == T_24222 ? T_23676_503 : GEN_2457;
  assign GEN_2459 = 9'h1f8 == T_24222 ? T_23676_504 : GEN_2458;
  assign GEN_2460 = 9'h1f9 == T_24222 ? T_23676_505 : GEN_2459;
  assign GEN_2461 = 9'h1fa == T_24222 ? T_23676_506 : GEN_2460;
  assign GEN_2462 = 9'h1fb == T_24222 ? T_23676_507 : GEN_2461;
  assign GEN_2463 = 9'h1fc == T_24222 ? T_23676_508 : GEN_2462;
  assign GEN_2464 = 9'h1fd == T_24222 ? T_23676_509 : GEN_2463;
  assign GEN_2465 = 9'h1fe == T_24222 ? T_23676_510 : GEN_2464;
  assign GEN_2466 = 9'h1ff == T_24222 ? T_23676_511 : GEN_2465;
  assign T_24260 = T_3205_bits_read ? GEN_5 : GEN_6;
  assign T_24261 = T_3205_ready & T_24257;
  assign T_24262 = T_3130_valid & T_24257;
  assign T_24263 = T_3169_ready & T_24260;
  assign T_24264 = T_3205_valid & T_24260;
  assign T_24266 = 512'h1 << T_24222;
  assign T_25293 = T_3130_valid & T_3205_ready;
  assign T_25294 = T_25293 & T_3205_bits_read;
  assign T_25295 = T_24266[0];
  assign T_25296 = T_25294 & T_25295;
  assign T_25299 = T_3205_bits_read == 1'h0;
  assign T_25300 = T_25293 & T_25299;
  assign T_25302 = T_25300 & T_25295;
  assign T_25303 = T_3205_valid & T_3169_ready;
  assign T_25304 = T_25303 & T_3205_bits_read;
  assign T_25306 = T_25304 & T_25295;
  assign T_25310 = T_25303 & T_25299;
  assign T_25312 = T_25310 & T_25295;
  assign T_25315 = T_24266[1];
  assign T_25316 = T_25294 & T_25315;
  assign T_25322 = T_25300 & T_25315;
  assign T_25326 = T_25304 & T_25315;
  assign T_25332 = T_25310 & T_25315;
  assign T_25335 = T_24266[2];
  assign T_25336 = T_25294 & T_25335;
  assign T_25342 = T_25300 & T_25335;
  assign T_25346 = T_25304 & T_25335;
  assign T_25352 = T_25310 & T_25335;
  assign T_25355 = T_24266[3];
  assign T_25356 = T_25294 & T_25355;
  assign T_25362 = T_25300 & T_25355;
  assign T_25366 = T_25304 & T_25355;
  assign T_25372 = T_25310 & T_25355;
  assign T_25375 = T_24266[4];
  assign T_25376 = T_25294 & T_25375;
  assign T_25382 = T_25300 & T_25375;
  assign T_25386 = T_25304 & T_25375;
  assign T_25392 = T_25310 & T_25375;
  assign T_25395 = T_24266[5];
  assign T_25396 = T_25294 & T_25395;
  assign T_25402 = T_25300 & T_25395;
  assign T_25406 = T_25304 & T_25395;
  assign T_25412 = T_25310 & T_25395;
  assign T_25415 = T_24266[6];
  assign T_25416 = T_25294 & T_25415;
  assign T_25422 = T_25300 & T_25415;
  assign T_25426 = T_25304 & T_25415;
  assign T_25432 = T_25310 & T_25415;
  assign T_25435 = T_24266[7];
  assign T_25436 = T_25294 & T_25435;
  assign T_25442 = T_25300 & T_25435;
  assign T_25446 = T_25304 & T_25435;
  assign T_25452 = T_25310 & T_25435;
  assign T_25455 = T_24266[8];
  assign T_25456 = T_25294 & T_25455;
  assign T_25462 = T_25300 & T_25455;
  assign T_25466 = T_25304 & T_25455;
  assign T_25472 = T_25310 & T_25455;
  assign T_25475 = T_24266[9];
  assign T_25476 = T_25294 & T_25475;
  assign T_25482 = T_25300 & T_25475;
  assign T_25486 = T_25304 & T_25475;
  assign T_25492 = T_25310 & T_25475;
  assign T_25495 = T_24266[10];
  assign T_25496 = T_25294 & T_25495;
  assign T_25502 = T_25300 & T_25495;
  assign T_25506 = T_25304 & T_25495;
  assign T_25512 = T_25310 & T_25495;
  assign T_25515 = T_24266[11];
  assign T_25516 = T_25294 & T_25515;
  assign T_25522 = T_25300 & T_25515;
  assign T_25526 = T_25304 & T_25515;
  assign T_25532 = T_25310 & T_25515;
  assign T_25535 = T_24266[12];
  assign T_25536 = T_25294 & T_25535;
  assign T_25542 = T_25300 & T_25535;
  assign T_25546 = T_25304 & T_25535;
  assign T_25552 = T_25310 & T_25535;
  assign T_25555 = T_24266[13];
  assign T_25556 = T_25294 & T_25555;
  assign T_25562 = T_25300 & T_25555;
  assign T_25566 = T_25304 & T_25555;
  assign T_25572 = T_25310 & T_25555;
  assign T_25575 = T_24266[14];
  assign T_25576 = T_25294 & T_25575;
  assign T_25582 = T_25300 & T_25575;
  assign T_25586 = T_25304 & T_25575;
  assign T_25592 = T_25310 & T_25575;
  assign T_25595 = T_24266[15];
  assign T_25596 = T_25294 & T_25595;
  assign T_25602 = T_25300 & T_25595;
  assign T_25606 = T_25304 & T_25595;
  assign T_25612 = T_25310 & T_25595;
  assign T_25615 = T_24266[16];
  assign T_25616 = T_25294 & T_25615;
  assign T_25622 = T_25300 & T_25615;
  assign T_25626 = T_25304 & T_25615;
  assign T_25632 = T_25310 & T_25615;
  assign T_25635 = T_24266[17];
  assign T_25636 = T_25294 & T_25635;
  assign T_25642 = T_25300 & T_25635;
  assign T_25646 = T_25304 & T_25635;
  assign T_25652 = T_25310 & T_25635;
  assign T_25655 = T_24266[18];
  assign T_25656 = T_25294 & T_25655;
  assign T_25662 = T_25300 & T_25655;
  assign T_25666 = T_25304 & T_25655;
  assign T_25672 = T_25310 & T_25655;
  assign T_25675 = T_24266[19];
  assign T_25676 = T_25294 & T_25675;
  assign T_25682 = T_25300 & T_25675;
  assign T_25686 = T_25304 & T_25675;
  assign T_25692 = T_25310 & T_25675;
  assign T_25695 = T_24266[20];
  assign T_25696 = T_25294 & T_25695;
  assign T_25702 = T_25300 & T_25695;
  assign T_25706 = T_25304 & T_25695;
  assign T_25712 = T_25310 & T_25695;
  assign T_25715 = T_24266[21];
  assign T_25716 = T_25294 & T_25715;
  assign T_25722 = T_25300 & T_25715;
  assign T_25726 = T_25304 & T_25715;
  assign T_25732 = T_25310 & T_25715;
  assign T_25735 = T_24266[22];
  assign T_25736 = T_25294 & T_25735;
  assign T_25742 = T_25300 & T_25735;
  assign T_25746 = T_25304 & T_25735;
  assign T_25752 = T_25310 & T_25735;
  assign T_25755 = T_24266[23];
  assign T_25756 = T_25294 & T_25755;
  assign T_25762 = T_25300 & T_25755;
  assign T_25766 = T_25304 & T_25755;
  assign T_25772 = T_25310 & T_25755;
  assign T_25775 = T_24266[24];
  assign T_25776 = T_25294 & T_25775;
  assign T_25782 = T_25300 & T_25775;
  assign T_25786 = T_25304 & T_25775;
  assign T_25792 = T_25310 & T_25775;
  assign T_25795 = T_24266[25];
  assign T_25796 = T_25294 & T_25795;
  assign T_25802 = T_25300 & T_25795;
  assign T_25806 = T_25304 & T_25795;
  assign T_25812 = T_25310 & T_25795;
  assign T_25815 = T_24266[26];
  assign T_25816 = T_25294 & T_25815;
  assign T_25822 = T_25300 & T_25815;
  assign T_25826 = T_25304 & T_25815;
  assign T_25832 = T_25310 & T_25815;
  assign T_25835 = T_24266[27];
  assign T_25836 = T_25294 & T_25835;
  assign T_25842 = T_25300 & T_25835;
  assign T_25846 = T_25304 & T_25835;
  assign T_25852 = T_25310 & T_25835;
  assign T_25855 = T_24266[28];
  assign T_25856 = T_25294 & T_25855;
  assign T_25862 = T_25300 & T_25855;
  assign T_25866 = T_25304 & T_25855;
  assign T_25872 = T_25310 & T_25855;
  assign T_25875 = T_24266[29];
  assign T_25876 = T_25294 & T_25875;
  assign T_25882 = T_25300 & T_25875;
  assign T_25886 = T_25304 & T_25875;
  assign T_25892 = T_25310 & T_25875;
  assign T_25895 = T_24266[30];
  assign T_25896 = T_25294 & T_25895;
  assign T_25902 = T_25300 & T_25895;
  assign T_25906 = T_25304 & T_25895;
  assign T_25912 = T_25310 & T_25895;
  assign T_25915 = T_24266[31];
  assign T_25916 = T_25294 & T_25915;
  assign T_25922 = T_25300 & T_25915;
  assign T_25926 = T_25304 & T_25915;
  assign T_25932 = T_25310 & T_25915;
  assign T_25935 = T_24266[32];
  assign T_25936 = T_25294 & T_25935;
  assign T_25942 = T_25300 & T_25935;
  assign T_25946 = T_25304 & T_25935;
  assign T_25952 = T_25310 & T_25935;
  assign T_25955 = T_24266[33];
  assign T_25956 = T_25294 & T_25955;
  assign T_25962 = T_25300 & T_25955;
  assign T_25966 = T_25304 & T_25955;
  assign T_25972 = T_25310 & T_25955;
  assign T_25975 = T_24266[34];
  assign T_25976 = T_25294 & T_25975;
  assign T_25982 = T_25300 & T_25975;
  assign T_25986 = T_25304 & T_25975;
  assign T_25992 = T_25310 & T_25975;
  assign T_25995 = T_24266[35];
  assign T_25996 = T_25294 & T_25995;
  assign T_26002 = T_25300 & T_25995;
  assign T_26006 = T_25304 & T_25995;
  assign T_26012 = T_25310 & T_25995;
  assign T_26015 = T_24266[36];
  assign T_26016 = T_25294 & T_26015;
  assign T_26022 = T_25300 & T_26015;
  assign T_26026 = T_25304 & T_26015;
  assign T_26032 = T_25310 & T_26015;
  assign T_26035 = T_24266[37];
  assign T_26036 = T_25294 & T_26035;
  assign T_26042 = T_25300 & T_26035;
  assign T_26046 = T_25304 & T_26035;
  assign T_26052 = T_25310 & T_26035;
  assign T_26055 = T_24266[38];
  assign T_26056 = T_25294 & T_26055;
  assign T_26062 = T_25300 & T_26055;
  assign T_26066 = T_25304 & T_26055;
  assign T_26072 = T_25310 & T_26055;
  assign T_26075 = T_24266[39];
  assign T_26076 = T_25294 & T_26075;
  assign T_26082 = T_25300 & T_26075;
  assign T_26086 = T_25304 & T_26075;
  assign T_26092 = T_25310 & T_26075;
  assign T_26095 = T_24266[40];
  assign T_26096 = T_25294 & T_26095;
  assign T_26102 = T_25300 & T_26095;
  assign T_26106 = T_25304 & T_26095;
  assign T_26112 = T_25310 & T_26095;
  assign T_26115 = T_24266[41];
  assign T_26116 = T_25294 & T_26115;
  assign T_26122 = T_25300 & T_26115;
  assign T_26126 = T_25304 & T_26115;
  assign T_26132 = T_25310 & T_26115;
  assign T_26135 = T_24266[42];
  assign T_26136 = T_25294 & T_26135;
  assign T_26142 = T_25300 & T_26135;
  assign T_26146 = T_25304 & T_26135;
  assign T_26152 = T_25310 & T_26135;
  assign T_26155 = T_24266[43];
  assign T_26156 = T_25294 & T_26155;
  assign T_26162 = T_25300 & T_26155;
  assign T_26166 = T_25304 & T_26155;
  assign T_26172 = T_25310 & T_26155;
  assign T_26175 = T_24266[44];
  assign T_26176 = T_25294 & T_26175;
  assign T_26182 = T_25300 & T_26175;
  assign T_26186 = T_25304 & T_26175;
  assign T_26192 = T_25310 & T_26175;
  assign T_26195 = T_24266[45];
  assign T_26196 = T_25294 & T_26195;
  assign T_26202 = T_25300 & T_26195;
  assign T_26206 = T_25304 & T_26195;
  assign T_26212 = T_25310 & T_26195;
  assign T_26215 = T_24266[46];
  assign T_26216 = T_25294 & T_26215;
  assign T_26222 = T_25300 & T_26215;
  assign T_26226 = T_25304 & T_26215;
  assign T_26232 = T_25310 & T_26215;
  assign T_26235 = T_24266[47];
  assign T_26236 = T_25294 & T_26235;
  assign T_26242 = T_25300 & T_26235;
  assign T_26246 = T_25304 & T_26235;
  assign T_26252 = T_25310 & T_26235;
  assign T_26255 = T_24266[48];
  assign T_26256 = T_25294 & T_26255;
  assign T_26262 = T_25300 & T_26255;
  assign T_26266 = T_25304 & T_26255;
  assign T_26272 = T_25310 & T_26255;
  assign T_26275 = T_24266[49];
  assign T_26276 = T_25294 & T_26275;
  assign T_26282 = T_25300 & T_26275;
  assign T_26286 = T_25304 & T_26275;
  assign T_26292 = T_25310 & T_26275;
  assign T_26295 = T_24266[50];
  assign T_26296 = T_25294 & T_26295;
  assign T_26302 = T_25300 & T_26295;
  assign T_26306 = T_25304 & T_26295;
  assign T_26312 = T_25310 & T_26295;
  assign T_26315 = T_24266[51];
  assign T_26316 = T_25294 & T_26315;
  assign T_26322 = T_25300 & T_26315;
  assign T_26326 = T_25304 & T_26315;
  assign T_26332 = T_25310 & T_26315;
  assign T_26575 = T_24266[64];
  assign T_26576 = T_25294 & T_26575;
  assign T_26582 = T_25300 & T_26575;
  assign T_26586 = T_25304 & T_26575;
  assign T_26592 = T_25310 & T_26575;
  assign T_26595 = T_24266[65];
  assign T_26596 = T_25294 & T_26595;
  assign T_26602 = T_25300 & T_26595;
  assign T_26606 = T_25304 & T_26595;
  assign T_26612 = T_25310 & T_26595;
  assign T_27855 = T_24266[128];
  assign T_27856 = T_25294 & T_27855;
  assign T_27862 = T_25300 & T_27855;
  assign T_27866 = T_25304 & T_27855;
  assign T_27872 = T_25310 & T_27855;
  assign T_27875 = T_24266[129];
  assign T_27876 = T_25294 & T_27875;
  assign T_27882 = T_25300 & T_27875;
  assign T_27886 = T_25304 & T_27875;
  assign T_27892 = T_25310 & T_27875;
  assign T_30415 = T_24266[256];
  assign T_30416 = T_25294 & T_30415;
  assign T_30422 = T_25300 & T_30415;
  assign T_30426 = T_25304 & T_30415;
  assign T_30432 = T_25310 & T_30415;
  assign T_30435 = T_24266[257];
  assign T_30436 = T_25294 & T_30435;
  assign T_30442 = T_25300 & T_30435;
  assign T_30446 = T_25304 & T_30435;
  assign T_30452 = T_25310 & T_30435;
  assign T_35533 = T_26576 & T_4319_31;
  assign T_35534 = T_35533 & T_4319_30;
  assign T_35535 = T_35534 & T_4319_29;
  assign T_35536 = T_35535 & T_4319_28;
  assign T_35537 = T_35536 & T_4319_27;
  assign T_35538 = T_35537 & T_4319_26;
  assign T_35539 = T_35538 & T_4319_25;
  assign T_35540 = T_35539 & T_4319_24;
  assign T_35541 = T_35540 & T_4319_23;
  assign T_35542 = T_35541 & T_4319_22;
  assign T_35543 = T_35542 & T_4319_21;
  assign T_35544 = T_35543 & T_4319_20;
  assign T_35545 = T_35544 & T_4319_19;
  assign T_35546 = T_35545 & T_4319_18;
  assign T_35547 = T_35546 & T_4319_17;
  assign T_35548 = T_35547 & T_4319_16;
  assign T_35549 = T_35548 & T_4319_15;
  assign T_35550 = T_35549 & T_4319_14;
  assign T_35551 = T_35550 & T_4319_13;
  assign T_35552 = T_35551 & T_4319_12;
  assign T_35553 = T_35552 & T_4319_11;
  assign T_35554 = T_35553 & T_4319_10;
  assign T_35555 = T_35554 & T_4319_9;
  assign T_35556 = T_35555 & T_4319_8;
  assign T_35557 = T_35556 & T_4319_7;
  assign T_35558 = T_35557 & T_4319_6;
  assign T_35559 = T_35558 & T_4319_5;
  assign T_35560 = T_35559 & T_4319_4;
  assign T_35561 = T_35560 & T_4319_3;
  assign T_35562 = T_35561 & T_4319_2;
  assign T_35563 = T_35562 & T_4319_1;
  assign T_35565 = T_26582 & T_4324_31;
  assign T_35566 = T_35565 & T_4324_30;
  assign T_35567 = T_35566 & T_4324_29;
  assign T_35568 = T_35567 & T_4324_28;
  assign T_35569 = T_35568 & T_4324_27;
  assign T_35570 = T_35569 & T_4324_26;
  assign T_35571 = T_35570 & T_4324_25;
  assign T_35572 = T_35571 & T_4324_24;
  assign T_35573 = T_35572 & T_4324_23;
  assign T_35574 = T_35573 & T_4324_22;
  assign T_35575 = T_35574 & T_4324_21;
  assign T_35576 = T_35575 & T_4324_20;
  assign T_35577 = T_35576 & T_4324_19;
  assign T_35578 = T_35577 & T_4324_18;
  assign T_35579 = T_35578 & T_4324_17;
  assign T_35580 = T_35579 & T_4324_16;
  assign T_35581 = T_35580 & T_4324_15;
  assign T_35582 = T_35581 & T_4324_14;
  assign T_35583 = T_35582 & T_4324_13;
  assign T_35584 = T_35583 & T_4324_12;
  assign T_35585 = T_35584 & T_4324_11;
  assign T_35586 = T_35585 & T_4324_10;
  assign T_35587 = T_35586 & T_4324_9;
  assign T_35588 = T_35587 & T_4324_8;
  assign T_35589 = T_35588 & T_4324_7;
  assign T_35590 = T_35589 & T_4324_6;
  assign T_35591 = T_35590 & T_4324_5;
  assign T_35592 = T_35591 & T_4324_4;
  assign T_35593 = T_35592 & T_4324_3;
  assign T_35594 = T_35593 & T_4324_2;
  assign T_35595 = T_35594 & T_4324_1;
  assign T_35597 = T_26586 & T_4329_31;
  assign T_35598 = T_35597 & T_4329_30;
  assign T_35599 = T_35598 & T_4329_29;
  assign T_35600 = T_35599 & T_4329_28;
  assign T_35601 = T_35600 & T_4329_27;
  assign T_35602 = T_35601 & T_4329_26;
  assign T_35603 = T_35602 & T_4329_25;
  assign T_35604 = T_35603 & T_4329_24;
  assign T_35605 = T_35604 & T_4329_23;
  assign T_35606 = T_35605 & T_4329_22;
  assign T_35607 = T_35606 & T_4329_21;
  assign T_35608 = T_35607 & T_4329_20;
  assign T_35609 = T_35608 & T_4329_19;
  assign T_35610 = T_35609 & T_4329_18;
  assign T_35611 = T_35610 & T_4329_17;
  assign T_35612 = T_35611 & T_4329_16;
  assign T_35613 = T_35612 & T_4329_15;
  assign T_35614 = T_35613 & T_4329_14;
  assign T_35615 = T_35614 & T_4329_13;
  assign T_35616 = T_35615 & T_4329_12;
  assign T_35617 = T_35616 & T_4329_11;
  assign T_35618 = T_35617 & T_4329_10;
  assign T_35619 = T_35618 & T_4329_9;
  assign T_35620 = T_35619 & T_4329_8;
  assign T_35621 = T_35620 & T_4329_7;
  assign T_35622 = T_35621 & T_4329_6;
  assign T_35623 = T_35622 & T_4329_5;
  assign T_35624 = T_35623 & T_4329_4;
  assign T_35625 = T_35624 & T_4329_3;
  assign T_35626 = T_35625 & T_4329_2;
  assign T_35627 = T_35626 & T_4329_1;
  assign T_35629 = T_26592 & T_4334_31;
  assign T_35630 = T_35629 & T_4334_30;
  assign T_35631 = T_35630 & T_4334_29;
  assign T_35632 = T_35631 & T_4334_28;
  assign T_35633 = T_35632 & T_4334_27;
  assign T_35634 = T_35633 & T_4334_26;
  assign T_35635 = T_35634 & T_4334_25;
  assign T_35636 = T_35635 & T_4334_24;
  assign T_35637 = T_35636 & T_4334_23;
  assign T_35638 = T_35637 & T_4334_22;
  assign T_35639 = T_35638 & T_4334_21;
  assign T_35640 = T_35639 & T_4334_20;
  assign T_35641 = T_35640 & T_4334_19;
  assign T_35642 = T_35641 & T_4334_18;
  assign T_35643 = T_35642 & T_4334_17;
  assign T_35644 = T_35643 & T_4334_16;
  assign T_35645 = T_35644 & T_4334_15;
  assign T_35646 = T_35645 & T_4334_14;
  assign T_35647 = T_35646 & T_4334_13;
  assign T_35648 = T_35647 & T_4334_12;
  assign T_35649 = T_35648 & T_4334_11;
  assign T_35650 = T_35649 & T_4334_10;
  assign T_35651 = T_35650 & T_4334_9;
  assign T_35652 = T_35651 & T_4334_8;
  assign T_35653 = T_35652 & T_4334_7;
  assign T_35654 = T_35653 & T_4334_6;
  assign T_35655 = T_35654 & T_4334_5;
  assign T_35656 = T_35655 & T_4334_4;
  assign T_35657 = T_35656 & T_4334_3;
  assign T_35658 = T_35657 & T_4334_2;
  assign T_35659 = T_35658 & T_4334_1;
  assign T_35691 = T_35562 & T_4319_0;
  assign T_35723 = T_35594 & T_4324_0;
  assign T_35755 = T_35626 & T_4329_0;
  assign T_35787 = T_35658 & T_4334_0;
  assign T_35818 = T_35561 & T_4319_1;
  assign T_35819 = T_35818 & T_4319_0;
  assign T_35850 = T_35593 & T_4324_1;
  assign T_35851 = T_35850 & T_4324_0;
  assign T_35882 = T_35625 & T_4329_1;
  assign T_35883 = T_35882 & T_4329_0;
  assign T_35914 = T_35657 & T_4334_1;
  assign T_35915 = T_35914 & T_4334_0;
  assign T_35945 = T_35560 & T_4319_2;
  assign T_35946 = T_35945 & T_4319_1;
  assign T_35947 = T_35946 & T_4319_0;
  assign T_35977 = T_35592 & T_4324_2;
  assign T_35978 = T_35977 & T_4324_1;
  assign T_35979 = T_35978 & T_4324_0;
  assign T_36009 = T_35624 & T_4329_2;
  assign T_36010 = T_36009 & T_4329_1;
  assign T_36011 = T_36010 & T_4329_0;
  assign T_36041 = T_35656 & T_4334_2;
  assign T_36042 = T_36041 & T_4334_1;
  assign T_36043 = T_36042 & T_4334_0;
  assign T_36072 = T_35559 & T_4319_3;
  assign T_36073 = T_36072 & T_4319_2;
  assign T_36074 = T_36073 & T_4319_1;
  assign T_36075 = T_36074 & T_4319_0;
  assign T_36104 = T_35591 & T_4324_3;
  assign T_36105 = T_36104 & T_4324_2;
  assign T_36106 = T_36105 & T_4324_1;
  assign T_36107 = T_36106 & T_4324_0;
  assign T_36136 = T_35623 & T_4329_3;
  assign T_36137 = T_36136 & T_4329_2;
  assign T_36138 = T_36137 & T_4329_1;
  assign T_36139 = T_36138 & T_4329_0;
  assign T_36168 = T_35655 & T_4334_3;
  assign T_36169 = T_36168 & T_4334_2;
  assign T_36170 = T_36169 & T_4334_1;
  assign T_36171 = T_36170 & T_4334_0;
  assign T_36199 = T_35558 & T_4319_4;
  assign T_36200 = T_36199 & T_4319_3;
  assign T_36201 = T_36200 & T_4319_2;
  assign T_36202 = T_36201 & T_4319_1;
  assign T_36203 = T_36202 & T_4319_0;
  assign T_36231 = T_35590 & T_4324_4;
  assign T_36232 = T_36231 & T_4324_3;
  assign T_36233 = T_36232 & T_4324_2;
  assign T_36234 = T_36233 & T_4324_1;
  assign T_36235 = T_36234 & T_4324_0;
  assign T_36263 = T_35622 & T_4329_4;
  assign T_36264 = T_36263 & T_4329_3;
  assign T_36265 = T_36264 & T_4329_2;
  assign T_36266 = T_36265 & T_4329_1;
  assign T_36267 = T_36266 & T_4329_0;
  assign T_36295 = T_35654 & T_4334_4;
  assign T_36296 = T_36295 & T_4334_3;
  assign T_36297 = T_36296 & T_4334_2;
  assign T_36298 = T_36297 & T_4334_1;
  assign T_36299 = T_36298 & T_4334_0;
  assign T_36326 = T_35557 & T_4319_5;
  assign T_36327 = T_36326 & T_4319_4;
  assign T_36328 = T_36327 & T_4319_3;
  assign T_36329 = T_36328 & T_4319_2;
  assign T_36330 = T_36329 & T_4319_1;
  assign T_36331 = T_36330 & T_4319_0;
  assign T_36358 = T_35589 & T_4324_5;
  assign T_36359 = T_36358 & T_4324_4;
  assign T_36360 = T_36359 & T_4324_3;
  assign T_36361 = T_36360 & T_4324_2;
  assign T_36362 = T_36361 & T_4324_1;
  assign T_36363 = T_36362 & T_4324_0;
  assign T_36390 = T_35621 & T_4329_5;
  assign T_36391 = T_36390 & T_4329_4;
  assign T_36392 = T_36391 & T_4329_3;
  assign T_36393 = T_36392 & T_4329_2;
  assign T_36394 = T_36393 & T_4329_1;
  assign T_36395 = T_36394 & T_4329_0;
  assign T_36422 = T_35653 & T_4334_5;
  assign T_36423 = T_36422 & T_4334_4;
  assign T_36424 = T_36423 & T_4334_3;
  assign T_36425 = T_36424 & T_4334_2;
  assign T_36426 = T_36425 & T_4334_1;
  assign T_36427 = T_36426 & T_4334_0;
  assign T_36453 = T_35556 & T_4319_6;
  assign T_36454 = T_36453 & T_4319_5;
  assign T_36455 = T_36454 & T_4319_4;
  assign T_36456 = T_36455 & T_4319_3;
  assign T_36457 = T_36456 & T_4319_2;
  assign T_36458 = T_36457 & T_4319_1;
  assign T_36459 = T_36458 & T_4319_0;
  assign T_36485 = T_35588 & T_4324_6;
  assign T_36486 = T_36485 & T_4324_5;
  assign T_36487 = T_36486 & T_4324_4;
  assign T_36488 = T_36487 & T_4324_3;
  assign T_36489 = T_36488 & T_4324_2;
  assign T_36490 = T_36489 & T_4324_1;
  assign T_36491 = T_36490 & T_4324_0;
  assign T_36517 = T_35620 & T_4329_6;
  assign T_36518 = T_36517 & T_4329_5;
  assign T_36519 = T_36518 & T_4329_4;
  assign T_36520 = T_36519 & T_4329_3;
  assign T_36521 = T_36520 & T_4329_2;
  assign T_36522 = T_36521 & T_4329_1;
  assign T_36523 = T_36522 & T_4329_0;
  assign T_36549 = T_35652 & T_4334_6;
  assign T_36550 = T_36549 & T_4334_5;
  assign T_36551 = T_36550 & T_4334_4;
  assign T_36552 = T_36551 & T_4334_3;
  assign T_36553 = T_36552 & T_4334_2;
  assign T_36554 = T_36553 & T_4334_1;
  assign T_36555 = T_36554 & T_4334_0;
  assign T_36580 = T_35555 & T_4319_7;
  assign T_36581 = T_36580 & T_4319_6;
  assign T_36582 = T_36581 & T_4319_5;
  assign T_36583 = T_36582 & T_4319_4;
  assign T_36584 = T_36583 & T_4319_3;
  assign T_36585 = T_36584 & T_4319_2;
  assign T_36586 = T_36585 & T_4319_1;
  assign T_36587 = T_36586 & T_4319_0;
  assign T_36612 = T_35587 & T_4324_7;
  assign T_36613 = T_36612 & T_4324_6;
  assign T_36614 = T_36613 & T_4324_5;
  assign T_36615 = T_36614 & T_4324_4;
  assign T_36616 = T_36615 & T_4324_3;
  assign T_36617 = T_36616 & T_4324_2;
  assign T_36618 = T_36617 & T_4324_1;
  assign T_36619 = T_36618 & T_4324_0;
  assign T_36644 = T_35619 & T_4329_7;
  assign T_36645 = T_36644 & T_4329_6;
  assign T_36646 = T_36645 & T_4329_5;
  assign T_36647 = T_36646 & T_4329_4;
  assign T_36648 = T_36647 & T_4329_3;
  assign T_36649 = T_36648 & T_4329_2;
  assign T_36650 = T_36649 & T_4329_1;
  assign T_36651 = T_36650 & T_4329_0;
  assign T_36676 = T_35651 & T_4334_7;
  assign T_36677 = T_36676 & T_4334_6;
  assign T_36678 = T_36677 & T_4334_5;
  assign T_36679 = T_36678 & T_4334_4;
  assign T_36680 = T_36679 & T_4334_3;
  assign T_36681 = T_36680 & T_4334_2;
  assign T_36682 = T_36681 & T_4334_1;
  assign T_36683 = T_36682 & T_4334_0;
  assign T_36707 = T_35554 & T_4319_8;
  assign T_36708 = T_36707 & T_4319_7;
  assign T_36709 = T_36708 & T_4319_6;
  assign T_36710 = T_36709 & T_4319_5;
  assign T_36711 = T_36710 & T_4319_4;
  assign T_36712 = T_36711 & T_4319_3;
  assign T_36713 = T_36712 & T_4319_2;
  assign T_36714 = T_36713 & T_4319_1;
  assign T_36715 = T_36714 & T_4319_0;
  assign T_36739 = T_35586 & T_4324_8;
  assign T_36740 = T_36739 & T_4324_7;
  assign T_36741 = T_36740 & T_4324_6;
  assign T_36742 = T_36741 & T_4324_5;
  assign T_36743 = T_36742 & T_4324_4;
  assign T_36744 = T_36743 & T_4324_3;
  assign T_36745 = T_36744 & T_4324_2;
  assign T_36746 = T_36745 & T_4324_1;
  assign T_36747 = T_36746 & T_4324_0;
  assign T_36771 = T_35618 & T_4329_8;
  assign T_36772 = T_36771 & T_4329_7;
  assign T_36773 = T_36772 & T_4329_6;
  assign T_36774 = T_36773 & T_4329_5;
  assign T_36775 = T_36774 & T_4329_4;
  assign T_36776 = T_36775 & T_4329_3;
  assign T_36777 = T_36776 & T_4329_2;
  assign T_36778 = T_36777 & T_4329_1;
  assign T_36779 = T_36778 & T_4329_0;
  assign T_36803 = T_35650 & T_4334_8;
  assign T_36804 = T_36803 & T_4334_7;
  assign T_36805 = T_36804 & T_4334_6;
  assign T_36806 = T_36805 & T_4334_5;
  assign T_36807 = T_36806 & T_4334_4;
  assign T_36808 = T_36807 & T_4334_3;
  assign T_36809 = T_36808 & T_4334_2;
  assign T_36810 = T_36809 & T_4334_1;
  assign T_36811 = T_36810 & T_4334_0;
  assign T_36834 = T_35553 & T_4319_9;
  assign T_36835 = T_36834 & T_4319_8;
  assign T_36836 = T_36835 & T_4319_7;
  assign T_36837 = T_36836 & T_4319_6;
  assign T_36838 = T_36837 & T_4319_5;
  assign T_36839 = T_36838 & T_4319_4;
  assign T_36840 = T_36839 & T_4319_3;
  assign T_36841 = T_36840 & T_4319_2;
  assign T_36842 = T_36841 & T_4319_1;
  assign T_36843 = T_36842 & T_4319_0;
  assign T_36866 = T_35585 & T_4324_9;
  assign T_36867 = T_36866 & T_4324_8;
  assign T_36868 = T_36867 & T_4324_7;
  assign T_36869 = T_36868 & T_4324_6;
  assign T_36870 = T_36869 & T_4324_5;
  assign T_36871 = T_36870 & T_4324_4;
  assign T_36872 = T_36871 & T_4324_3;
  assign T_36873 = T_36872 & T_4324_2;
  assign T_36874 = T_36873 & T_4324_1;
  assign T_36875 = T_36874 & T_4324_0;
  assign T_36898 = T_35617 & T_4329_9;
  assign T_36899 = T_36898 & T_4329_8;
  assign T_36900 = T_36899 & T_4329_7;
  assign T_36901 = T_36900 & T_4329_6;
  assign T_36902 = T_36901 & T_4329_5;
  assign T_36903 = T_36902 & T_4329_4;
  assign T_36904 = T_36903 & T_4329_3;
  assign T_36905 = T_36904 & T_4329_2;
  assign T_36906 = T_36905 & T_4329_1;
  assign T_36907 = T_36906 & T_4329_0;
  assign T_36930 = T_35649 & T_4334_9;
  assign T_36931 = T_36930 & T_4334_8;
  assign T_36932 = T_36931 & T_4334_7;
  assign T_36933 = T_36932 & T_4334_6;
  assign T_36934 = T_36933 & T_4334_5;
  assign T_36935 = T_36934 & T_4334_4;
  assign T_36936 = T_36935 & T_4334_3;
  assign T_36937 = T_36936 & T_4334_2;
  assign T_36938 = T_36937 & T_4334_1;
  assign T_36939 = T_36938 & T_4334_0;
  assign T_36961 = T_35552 & T_4319_10;
  assign T_36962 = T_36961 & T_4319_9;
  assign T_36963 = T_36962 & T_4319_8;
  assign T_36964 = T_36963 & T_4319_7;
  assign T_36965 = T_36964 & T_4319_6;
  assign T_36966 = T_36965 & T_4319_5;
  assign T_36967 = T_36966 & T_4319_4;
  assign T_36968 = T_36967 & T_4319_3;
  assign T_36969 = T_36968 & T_4319_2;
  assign T_36970 = T_36969 & T_4319_1;
  assign T_36971 = T_36970 & T_4319_0;
  assign T_36993 = T_35584 & T_4324_10;
  assign T_36994 = T_36993 & T_4324_9;
  assign T_36995 = T_36994 & T_4324_8;
  assign T_36996 = T_36995 & T_4324_7;
  assign T_36997 = T_36996 & T_4324_6;
  assign T_36998 = T_36997 & T_4324_5;
  assign T_36999 = T_36998 & T_4324_4;
  assign T_37000 = T_36999 & T_4324_3;
  assign T_37001 = T_37000 & T_4324_2;
  assign T_37002 = T_37001 & T_4324_1;
  assign T_37003 = T_37002 & T_4324_0;
  assign T_37025 = T_35616 & T_4329_10;
  assign T_37026 = T_37025 & T_4329_9;
  assign T_37027 = T_37026 & T_4329_8;
  assign T_37028 = T_37027 & T_4329_7;
  assign T_37029 = T_37028 & T_4329_6;
  assign T_37030 = T_37029 & T_4329_5;
  assign T_37031 = T_37030 & T_4329_4;
  assign T_37032 = T_37031 & T_4329_3;
  assign T_37033 = T_37032 & T_4329_2;
  assign T_37034 = T_37033 & T_4329_1;
  assign T_37035 = T_37034 & T_4329_0;
  assign T_37057 = T_35648 & T_4334_10;
  assign T_37058 = T_37057 & T_4334_9;
  assign T_37059 = T_37058 & T_4334_8;
  assign T_37060 = T_37059 & T_4334_7;
  assign T_37061 = T_37060 & T_4334_6;
  assign T_37062 = T_37061 & T_4334_5;
  assign T_37063 = T_37062 & T_4334_4;
  assign T_37064 = T_37063 & T_4334_3;
  assign T_37065 = T_37064 & T_4334_2;
  assign T_37066 = T_37065 & T_4334_1;
  assign T_37067 = T_37066 & T_4334_0;
  assign T_37088 = T_35551 & T_4319_11;
  assign T_37089 = T_37088 & T_4319_10;
  assign T_37090 = T_37089 & T_4319_9;
  assign T_37091 = T_37090 & T_4319_8;
  assign T_37092 = T_37091 & T_4319_7;
  assign T_37093 = T_37092 & T_4319_6;
  assign T_37094 = T_37093 & T_4319_5;
  assign T_37095 = T_37094 & T_4319_4;
  assign T_37096 = T_37095 & T_4319_3;
  assign T_37097 = T_37096 & T_4319_2;
  assign T_37098 = T_37097 & T_4319_1;
  assign T_37099 = T_37098 & T_4319_0;
  assign T_37120 = T_35583 & T_4324_11;
  assign T_37121 = T_37120 & T_4324_10;
  assign T_37122 = T_37121 & T_4324_9;
  assign T_37123 = T_37122 & T_4324_8;
  assign T_37124 = T_37123 & T_4324_7;
  assign T_37125 = T_37124 & T_4324_6;
  assign T_37126 = T_37125 & T_4324_5;
  assign T_37127 = T_37126 & T_4324_4;
  assign T_37128 = T_37127 & T_4324_3;
  assign T_37129 = T_37128 & T_4324_2;
  assign T_37130 = T_37129 & T_4324_1;
  assign T_37131 = T_37130 & T_4324_0;
  assign T_37152 = T_35615 & T_4329_11;
  assign T_37153 = T_37152 & T_4329_10;
  assign T_37154 = T_37153 & T_4329_9;
  assign T_37155 = T_37154 & T_4329_8;
  assign T_37156 = T_37155 & T_4329_7;
  assign T_37157 = T_37156 & T_4329_6;
  assign T_37158 = T_37157 & T_4329_5;
  assign T_37159 = T_37158 & T_4329_4;
  assign T_37160 = T_37159 & T_4329_3;
  assign T_37161 = T_37160 & T_4329_2;
  assign T_37162 = T_37161 & T_4329_1;
  assign T_37163 = T_37162 & T_4329_0;
  assign T_37184 = T_35647 & T_4334_11;
  assign T_37185 = T_37184 & T_4334_10;
  assign T_37186 = T_37185 & T_4334_9;
  assign T_37187 = T_37186 & T_4334_8;
  assign T_37188 = T_37187 & T_4334_7;
  assign T_37189 = T_37188 & T_4334_6;
  assign T_37190 = T_37189 & T_4334_5;
  assign T_37191 = T_37190 & T_4334_4;
  assign T_37192 = T_37191 & T_4334_3;
  assign T_37193 = T_37192 & T_4334_2;
  assign T_37194 = T_37193 & T_4334_1;
  assign T_37195 = T_37194 & T_4334_0;
  assign T_37215 = T_35550 & T_4319_12;
  assign T_37216 = T_37215 & T_4319_11;
  assign T_37217 = T_37216 & T_4319_10;
  assign T_37218 = T_37217 & T_4319_9;
  assign T_37219 = T_37218 & T_4319_8;
  assign T_37220 = T_37219 & T_4319_7;
  assign T_37221 = T_37220 & T_4319_6;
  assign T_37222 = T_37221 & T_4319_5;
  assign T_37223 = T_37222 & T_4319_4;
  assign T_37224 = T_37223 & T_4319_3;
  assign T_37225 = T_37224 & T_4319_2;
  assign T_37226 = T_37225 & T_4319_1;
  assign T_37227 = T_37226 & T_4319_0;
  assign T_37247 = T_35582 & T_4324_12;
  assign T_37248 = T_37247 & T_4324_11;
  assign T_37249 = T_37248 & T_4324_10;
  assign T_37250 = T_37249 & T_4324_9;
  assign T_37251 = T_37250 & T_4324_8;
  assign T_37252 = T_37251 & T_4324_7;
  assign T_37253 = T_37252 & T_4324_6;
  assign T_37254 = T_37253 & T_4324_5;
  assign T_37255 = T_37254 & T_4324_4;
  assign T_37256 = T_37255 & T_4324_3;
  assign T_37257 = T_37256 & T_4324_2;
  assign T_37258 = T_37257 & T_4324_1;
  assign T_37259 = T_37258 & T_4324_0;
  assign T_37279 = T_35614 & T_4329_12;
  assign T_37280 = T_37279 & T_4329_11;
  assign T_37281 = T_37280 & T_4329_10;
  assign T_37282 = T_37281 & T_4329_9;
  assign T_37283 = T_37282 & T_4329_8;
  assign T_37284 = T_37283 & T_4329_7;
  assign T_37285 = T_37284 & T_4329_6;
  assign T_37286 = T_37285 & T_4329_5;
  assign T_37287 = T_37286 & T_4329_4;
  assign T_37288 = T_37287 & T_4329_3;
  assign T_37289 = T_37288 & T_4329_2;
  assign T_37290 = T_37289 & T_4329_1;
  assign T_37291 = T_37290 & T_4329_0;
  assign T_37311 = T_35646 & T_4334_12;
  assign T_37312 = T_37311 & T_4334_11;
  assign T_37313 = T_37312 & T_4334_10;
  assign T_37314 = T_37313 & T_4334_9;
  assign T_37315 = T_37314 & T_4334_8;
  assign T_37316 = T_37315 & T_4334_7;
  assign T_37317 = T_37316 & T_4334_6;
  assign T_37318 = T_37317 & T_4334_5;
  assign T_37319 = T_37318 & T_4334_4;
  assign T_37320 = T_37319 & T_4334_3;
  assign T_37321 = T_37320 & T_4334_2;
  assign T_37322 = T_37321 & T_4334_1;
  assign T_37323 = T_37322 & T_4334_0;
  assign T_37342 = T_35549 & T_4319_13;
  assign T_37343 = T_37342 & T_4319_12;
  assign T_37344 = T_37343 & T_4319_11;
  assign T_37345 = T_37344 & T_4319_10;
  assign T_37346 = T_37345 & T_4319_9;
  assign T_37347 = T_37346 & T_4319_8;
  assign T_37348 = T_37347 & T_4319_7;
  assign T_37349 = T_37348 & T_4319_6;
  assign T_37350 = T_37349 & T_4319_5;
  assign T_37351 = T_37350 & T_4319_4;
  assign T_37352 = T_37351 & T_4319_3;
  assign T_37353 = T_37352 & T_4319_2;
  assign T_37354 = T_37353 & T_4319_1;
  assign T_37355 = T_37354 & T_4319_0;
  assign T_37374 = T_35581 & T_4324_13;
  assign T_37375 = T_37374 & T_4324_12;
  assign T_37376 = T_37375 & T_4324_11;
  assign T_37377 = T_37376 & T_4324_10;
  assign T_37378 = T_37377 & T_4324_9;
  assign T_37379 = T_37378 & T_4324_8;
  assign T_37380 = T_37379 & T_4324_7;
  assign T_37381 = T_37380 & T_4324_6;
  assign T_37382 = T_37381 & T_4324_5;
  assign T_37383 = T_37382 & T_4324_4;
  assign T_37384 = T_37383 & T_4324_3;
  assign T_37385 = T_37384 & T_4324_2;
  assign T_37386 = T_37385 & T_4324_1;
  assign T_37387 = T_37386 & T_4324_0;
  assign T_37406 = T_35613 & T_4329_13;
  assign T_37407 = T_37406 & T_4329_12;
  assign T_37408 = T_37407 & T_4329_11;
  assign T_37409 = T_37408 & T_4329_10;
  assign T_37410 = T_37409 & T_4329_9;
  assign T_37411 = T_37410 & T_4329_8;
  assign T_37412 = T_37411 & T_4329_7;
  assign T_37413 = T_37412 & T_4329_6;
  assign T_37414 = T_37413 & T_4329_5;
  assign T_37415 = T_37414 & T_4329_4;
  assign T_37416 = T_37415 & T_4329_3;
  assign T_37417 = T_37416 & T_4329_2;
  assign T_37418 = T_37417 & T_4329_1;
  assign T_37419 = T_37418 & T_4329_0;
  assign T_37438 = T_35645 & T_4334_13;
  assign T_37439 = T_37438 & T_4334_12;
  assign T_37440 = T_37439 & T_4334_11;
  assign T_37441 = T_37440 & T_4334_10;
  assign T_37442 = T_37441 & T_4334_9;
  assign T_37443 = T_37442 & T_4334_8;
  assign T_37444 = T_37443 & T_4334_7;
  assign T_37445 = T_37444 & T_4334_6;
  assign T_37446 = T_37445 & T_4334_5;
  assign T_37447 = T_37446 & T_4334_4;
  assign T_37448 = T_37447 & T_4334_3;
  assign T_37449 = T_37448 & T_4334_2;
  assign T_37450 = T_37449 & T_4334_1;
  assign T_37451 = T_37450 & T_4334_0;
  assign T_37469 = T_35548 & T_4319_14;
  assign T_37470 = T_37469 & T_4319_13;
  assign T_37471 = T_37470 & T_4319_12;
  assign T_37472 = T_37471 & T_4319_11;
  assign T_37473 = T_37472 & T_4319_10;
  assign T_37474 = T_37473 & T_4319_9;
  assign T_37475 = T_37474 & T_4319_8;
  assign T_37476 = T_37475 & T_4319_7;
  assign T_37477 = T_37476 & T_4319_6;
  assign T_37478 = T_37477 & T_4319_5;
  assign T_37479 = T_37478 & T_4319_4;
  assign T_37480 = T_37479 & T_4319_3;
  assign T_37481 = T_37480 & T_4319_2;
  assign T_37482 = T_37481 & T_4319_1;
  assign T_37483 = T_37482 & T_4319_0;
  assign T_37501 = T_35580 & T_4324_14;
  assign T_37502 = T_37501 & T_4324_13;
  assign T_37503 = T_37502 & T_4324_12;
  assign T_37504 = T_37503 & T_4324_11;
  assign T_37505 = T_37504 & T_4324_10;
  assign T_37506 = T_37505 & T_4324_9;
  assign T_37507 = T_37506 & T_4324_8;
  assign T_37508 = T_37507 & T_4324_7;
  assign T_37509 = T_37508 & T_4324_6;
  assign T_37510 = T_37509 & T_4324_5;
  assign T_37511 = T_37510 & T_4324_4;
  assign T_37512 = T_37511 & T_4324_3;
  assign T_37513 = T_37512 & T_4324_2;
  assign T_37514 = T_37513 & T_4324_1;
  assign T_37515 = T_37514 & T_4324_0;
  assign T_37533 = T_35612 & T_4329_14;
  assign T_37534 = T_37533 & T_4329_13;
  assign T_37535 = T_37534 & T_4329_12;
  assign T_37536 = T_37535 & T_4329_11;
  assign T_37537 = T_37536 & T_4329_10;
  assign T_37538 = T_37537 & T_4329_9;
  assign T_37539 = T_37538 & T_4329_8;
  assign T_37540 = T_37539 & T_4329_7;
  assign T_37541 = T_37540 & T_4329_6;
  assign T_37542 = T_37541 & T_4329_5;
  assign T_37543 = T_37542 & T_4329_4;
  assign T_37544 = T_37543 & T_4329_3;
  assign T_37545 = T_37544 & T_4329_2;
  assign T_37546 = T_37545 & T_4329_1;
  assign T_37547 = T_37546 & T_4329_0;
  assign T_37565 = T_35644 & T_4334_14;
  assign T_37566 = T_37565 & T_4334_13;
  assign T_37567 = T_37566 & T_4334_12;
  assign T_37568 = T_37567 & T_4334_11;
  assign T_37569 = T_37568 & T_4334_10;
  assign T_37570 = T_37569 & T_4334_9;
  assign T_37571 = T_37570 & T_4334_8;
  assign T_37572 = T_37571 & T_4334_7;
  assign T_37573 = T_37572 & T_4334_6;
  assign T_37574 = T_37573 & T_4334_5;
  assign T_37575 = T_37574 & T_4334_4;
  assign T_37576 = T_37575 & T_4334_3;
  assign T_37577 = T_37576 & T_4334_2;
  assign T_37578 = T_37577 & T_4334_1;
  assign T_37579 = T_37578 & T_4334_0;
  assign T_37596 = T_35547 & T_4319_15;
  assign T_37597 = T_37596 & T_4319_14;
  assign T_37598 = T_37597 & T_4319_13;
  assign T_37599 = T_37598 & T_4319_12;
  assign T_37600 = T_37599 & T_4319_11;
  assign T_37601 = T_37600 & T_4319_10;
  assign T_37602 = T_37601 & T_4319_9;
  assign T_37603 = T_37602 & T_4319_8;
  assign T_37604 = T_37603 & T_4319_7;
  assign T_37605 = T_37604 & T_4319_6;
  assign T_37606 = T_37605 & T_4319_5;
  assign T_37607 = T_37606 & T_4319_4;
  assign T_37608 = T_37607 & T_4319_3;
  assign T_37609 = T_37608 & T_4319_2;
  assign T_37610 = T_37609 & T_4319_1;
  assign T_37611 = T_37610 & T_4319_0;
  assign T_37628 = T_35579 & T_4324_15;
  assign T_37629 = T_37628 & T_4324_14;
  assign T_37630 = T_37629 & T_4324_13;
  assign T_37631 = T_37630 & T_4324_12;
  assign T_37632 = T_37631 & T_4324_11;
  assign T_37633 = T_37632 & T_4324_10;
  assign T_37634 = T_37633 & T_4324_9;
  assign T_37635 = T_37634 & T_4324_8;
  assign T_37636 = T_37635 & T_4324_7;
  assign T_37637 = T_37636 & T_4324_6;
  assign T_37638 = T_37637 & T_4324_5;
  assign T_37639 = T_37638 & T_4324_4;
  assign T_37640 = T_37639 & T_4324_3;
  assign T_37641 = T_37640 & T_4324_2;
  assign T_37642 = T_37641 & T_4324_1;
  assign T_37643 = T_37642 & T_4324_0;
  assign T_37660 = T_35611 & T_4329_15;
  assign T_37661 = T_37660 & T_4329_14;
  assign T_37662 = T_37661 & T_4329_13;
  assign T_37663 = T_37662 & T_4329_12;
  assign T_37664 = T_37663 & T_4329_11;
  assign T_37665 = T_37664 & T_4329_10;
  assign T_37666 = T_37665 & T_4329_9;
  assign T_37667 = T_37666 & T_4329_8;
  assign T_37668 = T_37667 & T_4329_7;
  assign T_37669 = T_37668 & T_4329_6;
  assign T_37670 = T_37669 & T_4329_5;
  assign T_37671 = T_37670 & T_4329_4;
  assign T_37672 = T_37671 & T_4329_3;
  assign T_37673 = T_37672 & T_4329_2;
  assign T_37674 = T_37673 & T_4329_1;
  assign T_37675 = T_37674 & T_4329_0;
  assign T_37692 = T_35643 & T_4334_15;
  assign T_37693 = T_37692 & T_4334_14;
  assign T_37694 = T_37693 & T_4334_13;
  assign T_37695 = T_37694 & T_4334_12;
  assign T_37696 = T_37695 & T_4334_11;
  assign T_37697 = T_37696 & T_4334_10;
  assign T_37698 = T_37697 & T_4334_9;
  assign T_37699 = T_37698 & T_4334_8;
  assign T_37700 = T_37699 & T_4334_7;
  assign T_37701 = T_37700 & T_4334_6;
  assign T_37702 = T_37701 & T_4334_5;
  assign T_37703 = T_37702 & T_4334_4;
  assign T_37704 = T_37703 & T_4334_3;
  assign T_37705 = T_37704 & T_4334_2;
  assign T_37706 = T_37705 & T_4334_1;
  assign T_37707 = T_37706 & T_4334_0;
  assign T_37723 = T_35546 & T_4319_16;
  assign T_37724 = T_37723 & T_4319_15;
  assign T_37725 = T_37724 & T_4319_14;
  assign T_37726 = T_37725 & T_4319_13;
  assign T_37727 = T_37726 & T_4319_12;
  assign T_37728 = T_37727 & T_4319_11;
  assign T_37729 = T_37728 & T_4319_10;
  assign T_37730 = T_37729 & T_4319_9;
  assign T_37731 = T_37730 & T_4319_8;
  assign T_37732 = T_37731 & T_4319_7;
  assign T_37733 = T_37732 & T_4319_6;
  assign T_37734 = T_37733 & T_4319_5;
  assign T_37735 = T_37734 & T_4319_4;
  assign T_37736 = T_37735 & T_4319_3;
  assign T_37737 = T_37736 & T_4319_2;
  assign T_37738 = T_37737 & T_4319_1;
  assign T_37739 = T_37738 & T_4319_0;
  assign T_37755 = T_35578 & T_4324_16;
  assign T_37756 = T_37755 & T_4324_15;
  assign T_37757 = T_37756 & T_4324_14;
  assign T_37758 = T_37757 & T_4324_13;
  assign T_37759 = T_37758 & T_4324_12;
  assign T_37760 = T_37759 & T_4324_11;
  assign T_37761 = T_37760 & T_4324_10;
  assign T_37762 = T_37761 & T_4324_9;
  assign T_37763 = T_37762 & T_4324_8;
  assign T_37764 = T_37763 & T_4324_7;
  assign T_37765 = T_37764 & T_4324_6;
  assign T_37766 = T_37765 & T_4324_5;
  assign T_37767 = T_37766 & T_4324_4;
  assign T_37768 = T_37767 & T_4324_3;
  assign T_37769 = T_37768 & T_4324_2;
  assign T_37770 = T_37769 & T_4324_1;
  assign T_37771 = T_37770 & T_4324_0;
  assign T_37787 = T_35610 & T_4329_16;
  assign T_37788 = T_37787 & T_4329_15;
  assign T_37789 = T_37788 & T_4329_14;
  assign T_37790 = T_37789 & T_4329_13;
  assign T_37791 = T_37790 & T_4329_12;
  assign T_37792 = T_37791 & T_4329_11;
  assign T_37793 = T_37792 & T_4329_10;
  assign T_37794 = T_37793 & T_4329_9;
  assign T_37795 = T_37794 & T_4329_8;
  assign T_37796 = T_37795 & T_4329_7;
  assign T_37797 = T_37796 & T_4329_6;
  assign T_37798 = T_37797 & T_4329_5;
  assign T_37799 = T_37798 & T_4329_4;
  assign T_37800 = T_37799 & T_4329_3;
  assign T_37801 = T_37800 & T_4329_2;
  assign T_37802 = T_37801 & T_4329_1;
  assign T_37803 = T_37802 & T_4329_0;
  assign T_37819 = T_35642 & T_4334_16;
  assign T_37820 = T_37819 & T_4334_15;
  assign T_37821 = T_37820 & T_4334_14;
  assign T_37822 = T_37821 & T_4334_13;
  assign T_37823 = T_37822 & T_4334_12;
  assign T_37824 = T_37823 & T_4334_11;
  assign T_37825 = T_37824 & T_4334_10;
  assign T_37826 = T_37825 & T_4334_9;
  assign T_37827 = T_37826 & T_4334_8;
  assign T_37828 = T_37827 & T_4334_7;
  assign T_37829 = T_37828 & T_4334_6;
  assign T_37830 = T_37829 & T_4334_5;
  assign T_37831 = T_37830 & T_4334_4;
  assign T_37832 = T_37831 & T_4334_3;
  assign T_37833 = T_37832 & T_4334_2;
  assign T_37834 = T_37833 & T_4334_1;
  assign T_37835 = T_37834 & T_4334_0;
  assign T_37850 = T_35545 & T_4319_17;
  assign T_37851 = T_37850 & T_4319_16;
  assign T_37852 = T_37851 & T_4319_15;
  assign T_37853 = T_37852 & T_4319_14;
  assign T_37854 = T_37853 & T_4319_13;
  assign T_37855 = T_37854 & T_4319_12;
  assign T_37856 = T_37855 & T_4319_11;
  assign T_37857 = T_37856 & T_4319_10;
  assign T_37858 = T_37857 & T_4319_9;
  assign T_37859 = T_37858 & T_4319_8;
  assign T_37860 = T_37859 & T_4319_7;
  assign T_37861 = T_37860 & T_4319_6;
  assign T_37862 = T_37861 & T_4319_5;
  assign T_37863 = T_37862 & T_4319_4;
  assign T_37864 = T_37863 & T_4319_3;
  assign T_37865 = T_37864 & T_4319_2;
  assign T_37866 = T_37865 & T_4319_1;
  assign T_37867 = T_37866 & T_4319_0;
  assign T_37882 = T_35577 & T_4324_17;
  assign T_37883 = T_37882 & T_4324_16;
  assign T_37884 = T_37883 & T_4324_15;
  assign T_37885 = T_37884 & T_4324_14;
  assign T_37886 = T_37885 & T_4324_13;
  assign T_37887 = T_37886 & T_4324_12;
  assign T_37888 = T_37887 & T_4324_11;
  assign T_37889 = T_37888 & T_4324_10;
  assign T_37890 = T_37889 & T_4324_9;
  assign T_37891 = T_37890 & T_4324_8;
  assign T_37892 = T_37891 & T_4324_7;
  assign T_37893 = T_37892 & T_4324_6;
  assign T_37894 = T_37893 & T_4324_5;
  assign T_37895 = T_37894 & T_4324_4;
  assign T_37896 = T_37895 & T_4324_3;
  assign T_37897 = T_37896 & T_4324_2;
  assign T_37898 = T_37897 & T_4324_1;
  assign T_37899 = T_37898 & T_4324_0;
  assign T_37914 = T_35609 & T_4329_17;
  assign T_37915 = T_37914 & T_4329_16;
  assign T_37916 = T_37915 & T_4329_15;
  assign T_37917 = T_37916 & T_4329_14;
  assign T_37918 = T_37917 & T_4329_13;
  assign T_37919 = T_37918 & T_4329_12;
  assign T_37920 = T_37919 & T_4329_11;
  assign T_37921 = T_37920 & T_4329_10;
  assign T_37922 = T_37921 & T_4329_9;
  assign T_37923 = T_37922 & T_4329_8;
  assign T_37924 = T_37923 & T_4329_7;
  assign T_37925 = T_37924 & T_4329_6;
  assign T_37926 = T_37925 & T_4329_5;
  assign T_37927 = T_37926 & T_4329_4;
  assign T_37928 = T_37927 & T_4329_3;
  assign T_37929 = T_37928 & T_4329_2;
  assign T_37930 = T_37929 & T_4329_1;
  assign T_37931 = T_37930 & T_4329_0;
  assign T_37946 = T_35641 & T_4334_17;
  assign T_37947 = T_37946 & T_4334_16;
  assign T_37948 = T_37947 & T_4334_15;
  assign T_37949 = T_37948 & T_4334_14;
  assign T_37950 = T_37949 & T_4334_13;
  assign T_37951 = T_37950 & T_4334_12;
  assign T_37952 = T_37951 & T_4334_11;
  assign T_37953 = T_37952 & T_4334_10;
  assign T_37954 = T_37953 & T_4334_9;
  assign T_37955 = T_37954 & T_4334_8;
  assign T_37956 = T_37955 & T_4334_7;
  assign T_37957 = T_37956 & T_4334_6;
  assign T_37958 = T_37957 & T_4334_5;
  assign T_37959 = T_37958 & T_4334_4;
  assign T_37960 = T_37959 & T_4334_3;
  assign T_37961 = T_37960 & T_4334_2;
  assign T_37962 = T_37961 & T_4334_1;
  assign T_37963 = T_37962 & T_4334_0;
  assign T_37977 = T_35544 & T_4319_18;
  assign T_37978 = T_37977 & T_4319_17;
  assign T_37979 = T_37978 & T_4319_16;
  assign T_37980 = T_37979 & T_4319_15;
  assign T_37981 = T_37980 & T_4319_14;
  assign T_37982 = T_37981 & T_4319_13;
  assign T_37983 = T_37982 & T_4319_12;
  assign T_37984 = T_37983 & T_4319_11;
  assign T_37985 = T_37984 & T_4319_10;
  assign T_37986 = T_37985 & T_4319_9;
  assign T_37987 = T_37986 & T_4319_8;
  assign T_37988 = T_37987 & T_4319_7;
  assign T_37989 = T_37988 & T_4319_6;
  assign T_37990 = T_37989 & T_4319_5;
  assign T_37991 = T_37990 & T_4319_4;
  assign T_37992 = T_37991 & T_4319_3;
  assign T_37993 = T_37992 & T_4319_2;
  assign T_37994 = T_37993 & T_4319_1;
  assign T_37995 = T_37994 & T_4319_0;
  assign T_38009 = T_35576 & T_4324_18;
  assign T_38010 = T_38009 & T_4324_17;
  assign T_38011 = T_38010 & T_4324_16;
  assign T_38012 = T_38011 & T_4324_15;
  assign T_38013 = T_38012 & T_4324_14;
  assign T_38014 = T_38013 & T_4324_13;
  assign T_38015 = T_38014 & T_4324_12;
  assign T_38016 = T_38015 & T_4324_11;
  assign T_38017 = T_38016 & T_4324_10;
  assign T_38018 = T_38017 & T_4324_9;
  assign T_38019 = T_38018 & T_4324_8;
  assign T_38020 = T_38019 & T_4324_7;
  assign T_38021 = T_38020 & T_4324_6;
  assign T_38022 = T_38021 & T_4324_5;
  assign T_38023 = T_38022 & T_4324_4;
  assign T_38024 = T_38023 & T_4324_3;
  assign T_38025 = T_38024 & T_4324_2;
  assign T_38026 = T_38025 & T_4324_1;
  assign T_38027 = T_38026 & T_4324_0;
  assign T_38041 = T_35608 & T_4329_18;
  assign T_38042 = T_38041 & T_4329_17;
  assign T_38043 = T_38042 & T_4329_16;
  assign T_38044 = T_38043 & T_4329_15;
  assign T_38045 = T_38044 & T_4329_14;
  assign T_38046 = T_38045 & T_4329_13;
  assign T_38047 = T_38046 & T_4329_12;
  assign T_38048 = T_38047 & T_4329_11;
  assign T_38049 = T_38048 & T_4329_10;
  assign T_38050 = T_38049 & T_4329_9;
  assign T_38051 = T_38050 & T_4329_8;
  assign T_38052 = T_38051 & T_4329_7;
  assign T_38053 = T_38052 & T_4329_6;
  assign T_38054 = T_38053 & T_4329_5;
  assign T_38055 = T_38054 & T_4329_4;
  assign T_38056 = T_38055 & T_4329_3;
  assign T_38057 = T_38056 & T_4329_2;
  assign T_38058 = T_38057 & T_4329_1;
  assign T_38059 = T_38058 & T_4329_0;
  assign T_38073 = T_35640 & T_4334_18;
  assign T_38074 = T_38073 & T_4334_17;
  assign T_38075 = T_38074 & T_4334_16;
  assign T_38076 = T_38075 & T_4334_15;
  assign T_38077 = T_38076 & T_4334_14;
  assign T_38078 = T_38077 & T_4334_13;
  assign T_38079 = T_38078 & T_4334_12;
  assign T_38080 = T_38079 & T_4334_11;
  assign T_38081 = T_38080 & T_4334_10;
  assign T_38082 = T_38081 & T_4334_9;
  assign T_38083 = T_38082 & T_4334_8;
  assign T_38084 = T_38083 & T_4334_7;
  assign T_38085 = T_38084 & T_4334_6;
  assign T_38086 = T_38085 & T_4334_5;
  assign T_38087 = T_38086 & T_4334_4;
  assign T_38088 = T_38087 & T_4334_3;
  assign T_38089 = T_38088 & T_4334_2;
  assign T_38090 = T_38089 & T_4334_1;
  assign T_38091 = T_38090 & T_4334_0;
  assign T_38104 = T_35543 & T_4319_19;
  assign T_38105 = T_38104 & T_4319_18;
  assign T_38106 = T_38105 & T_4319_17;
  assign T_38107 = T_38106 & T_4319_16;
  assign T_38108 = T_38107 & T_4319_15;
  assign T_38109 = T_38108 & T_4319_14;
  assign T_38110 = T_38109 & T_4319_13;
  assign T_38111 = T_38110 & T_4319_12;
  assign T_38112 = T_38111 & T_4319_11;
  assign T_38113 = T_38112 & T_4319_10;
  assign T_38114 = T_38113 & T_4319_9;
  assign T_38115 = T_38114 & T_4319_8;
  assign T_38116 = T_38115 & T_4319_7;
  assign T_38117 = T_38116 & T_4319_6;
  assign T_38118 = T_38117 & T_4319_5;
  assign T_38119 = T_38118 & T_4319_4;
  assign T_38120 = T_38119 & T_4319_3;
  assign T_38121 = T_38120 & T_4319_2;
  assign T_38122 = T_38121 & T_4319_1;
  assign T_38123 = T_38122 & T_4319_0;
  assign T_38136 = T_35575 & T_4324_19;
  assign T_38137 = T_38136 & T_4324_18;
  assign T_38138 = T_38137 & T_4324_17;
  assign T_38139 = T_38138 & T_4324_16;
  assign T_38140 = T_38139 & T_4324_15;
  assign T_38141 = T_38140 & T_4324_14;
  assign T_38142 = T_38141 & T_4324_13;
  assign T_38143 = T_38142 & T_4324_12;
  assign T_38144 = T_38143 & T_4324_11;
  assign T_38145 = T_38144 & T_4324_10;
  assign T_38146 = T_38145 & T_4324_9;
  assign T_38147 = T_38146 & T_4324_8;
  assign T_38148 = T_38147 & T_4324_7;
  assign T_38149 = T_38148 & T_4324_6;
  assign T_38150 = T_38149 & T_4324_5;
  assign T_38151 = T_38150 & T_4324_4;
  assign T_38152 = T_38151 & T_4324_3;
  assign T_38153 = T_38152 & T_4324_2;
  assign T_38154 = T_38153 & T_4324_1;
  assign T_38155 = T_38154 & T_4324_0;
  assign T_38168 = T_35607 & T_4329_19;
  assign T_38169 = T_38168 & T_4329_18;
  assign T_38170 = T_38169 & T_4329_17;
  assign T_38171 = T_38170 & T_4329_16;
  assign T_38172 = T_38171 & T_4329_15;
  assign T_38173 = T_38172 & T_4329_14;
  assign T_38174 = T_38173 & T_4329_13;
  assign T_38175 = T_38174 & T_4329_12;
  assign T_38176 = T_38175 & T_4329_11;
  assign T_38177 = T_38176 & T_4329_10;
  assign T_38178 = T_38177 & T_4329_9;
  assign T_38179 = T_38178 & T_4329_8;
  assign T_38180 = T_38179 & T_4329_7;
  assign T_38181 = T_38180 & T_4329_6;
  assign T_38182 = T_38181 & T_4329_5;
  assign T_38183 = T_38182 & T_4329_4;
  assign T_38184 = T_38183 & T_4329_3;
  assign T_38185 = T_38184 & T_4329_2;
  assign T_38186 = T_38185 & T_4329_1;
  assign T_38187 = T_38186 & T_4329_0;
  assign T_38200 = T_35639 & T_4334_19;
  assign T_38201 = T_38200 & T_4334_18;
  assign T_38202 = T_38201 & T_4334_17;
  assign T_38203 = T_38202 & T_4334_16;
  assign T_38204 = T_38203 & T_4334_15;
  assign T_38205 = T_38204 & T_4334_14;
  assign T_38206 = T_38205 & T_4334_13;
  assign T_38207 = T_38206 & T_4334_12;
  assign T_38208 = T_38207 & T_4334_11;
  assign T_38209 = T_38208 & T_4334_10;
  assign T_38210 = T_38209 & T_4334_9;
  assign T_38211 = T_38210 & T_4334_8;
  assign T_38212 = T_38211 & T_4334_7;
  assign T_38213 = T_38212 & T_4334_6;
  assign T_38214 = T_38213 & T_4334_5;
  assign T_38215 = T_38214 & T_4334_4;
  assign T_38216 = T_38215 & T_4334_3;
  assign T_38217 = T_38216 & T_4334_2;
  assign T_38218 = T_38217 & T_4334_1;
  assign T_38219 = T_38218 & T_4334_0;
  assign T_38231 = T_35542 & T_4319_20;
  assign T_38232 = T_38231 & T_4319_19;
  assign T_38233 = T_38232 & T_4319_18;
  assign T_38234 = T_38233 & T_4319_17;
  assign T_38235 = T_38234 & T_4319_16;
  assign T_38236 = T_38235 & T_4319_15;
  assign T_38237 = T_38236 & T_4319_14;
  assign T_38238 = T_38237 & T_4319_13;
  assign T_38239 = T_38238 & T_4319_12;
  assign T_38240 = T_38239 & T_4319_11;
  assign T_38241 = T_38240 & T_4319_10;
  assign T_38242 = T_38241 & T_4319_9;
  assign T_38243 = T_38242 & T_4319_8;
  assign T_38244 = T_38243 & T_4319_7;
  assign T_38245 = T_38244 & T_4319_6;
  assign T_38246 = T_38245 & T_4319_5;
  assign T_38247 = T_38246 & T_4319_4;
  assign T_38248 = T_38247 & T_4319_3;
  assign T_38249 = T_38248 & T_4319_2;
  assign T_38250 = T_38249 & T_4319_1;
  assign T_38251 = T_38250 & T_4319_0;
  assign T_38263 = T_35574 & T_4324_20;
  assign T_38264 = T_38263 & T_4324_19;
  assign T_38265 = T_38264 & T_4324_18;
  assign T_38266 = T_38265 & T_4324_17;
  assign T_38267 = T_38266 & T_4324_16;
  assign T_38268 = T_38267 & T_4324_15;
  assign T_38269 = T_38268 & T_4324_14;
  assign T_38270 = T_38269 & T_4324_13;
  assign T_38271 = T_38270 & T_4324_12;
  assign T_38272 = T_38271 & T_4324_11;
  assign T_38273 = T_38272 & T_4324_10;
  assign T_38274 = T_38273 & T_4324_9;
  assign T_38275 = T_38274 & T_4324_8;
  assign T_38276 = T_38275 & T_4324_7;
  assign T_38277 = T_38276 & T_4324_6;
  assign T_38278 = T_38277 & T_4324_5;
  assign T_38279 = T_38278 & T_4324_4;
  assign T_38280 = T_38279 & T_4324_3;
  assign T_38281 = T_38280 & T_4324_2;
  assign T_38282 = T_38281 & T_4324_1;
  assign T_38283 = T_38282 & T_4324_0;
  assign T_38295 = T_35606 & T_4329_20;
  assign T_38296 = T_38295 & T_4329_19;
  assign T_38297 = T_38296 & T_4329_18;
  assign T_38298 = T_38297 & T_4329_17;
  assign T_38299 = T_38298 & T_4329_16;
  assign T_38300 = T_38299 & T_4329_15;
  assign T_38301 = T_38300 & T_4329_14;
  assign T_38302 = T_38301 & T_4329_13;
  assign T_38303 = T_38302 & T_4329_12;
  assign T_38304 = T_38303 & T_4329_11;
  assign T_38305 = T_38304 & T_4329_10;
  assign T_38306 = T_38305 & T_4329_9;
  assign T_38307 = T_38306 & T_4329_8;
  assign T_38308 = T_38307 & T_4329_7;
  assign T_38309 = T_38308 & T_4329_6;
  assign T_38310 = T_38309 & T_4329_5;
  assign T_38311 = T_38310 & T_4329_4;
  assign T_38312 = T_38311 & T_4329_3;
  assign T_38313 = T_38312 & T_4329_2;
  assign T_38314 = T_38313 & T_4329_1;
  assign T_38315 = T_38314 & T_4329_0;
  assign T_38327 = T_35638 & T_4334_20;
  assign T_38328 = T_38327 & T_4334_19;
  assign T_38329 = T_38328 & T_4334_18;
  assign T_38330 = T_38329 & T_4334_17;
  assign T_38331 = T_38330 & T_4334_16;
  assign T_38332 = T_38331 & T_4334_15;
  assign T_38333 = T_38332 & T_4334_14;
  assign T_38334 = T_38333 & T_4334_13;
  assign T_38335 = T_38334 & T_4334_12;
  assign T_38336 = T_38335 & T_4334_11;
  assign T_38337 = T_38336 & T_4334_10;
  assign T_38338 = T_38337 & T_4334_9;
  assign T_38339 = T_38338 & T_4334_8;
  assign T_38340 = T_38339 & T_4334_7;
  assign T_38341 = T_38340 & T_4334_6;
  assign T_38342 = T_38341 & T_4334_5;
  assign T_38343 = T_38342 & T_4334_4;
  assign T_38344 = T_38343 & T_4334_3;
  assign T_38345 = T_38344 & T_4334_2;
  assign T_38346 = T_38345 & T_4334_1;
  assign T_38347 = T_38346 & T_4334_0;
  assign T_38358 = T_35541 & T_4319_21;
  assign T_38359 = T_38358 & T_4319_20;
  assign T_38360 = T_38359 & T_4319_19;
  assign T_38361 = T_38360 & T_4319_18;
  assign T_38362 = T_38361 & T_4319_17;
  assign T_38363 = T_38362 & T_4319_16;
  assign T_38364 = T_38363 & T_4319_15;
  assign T_38365 = T_38364 & T_4319_14;
  assign T_38366 = T_38365 & T_4319_13;
  assign T_38367 = T_38366 & T_4319_12;
  assign T_38368 = T_38367 & T_4319_11;
  assign T_38369 = T_38368 & T_4319_10;
  assign T_38370 = T_38369 & T_4319_9;
  assign T_38371 = T_38370 & T_4319_8;
  assign T_38372 = T_38371 & T_4319_7;
  assign T_38373 = T_38372 & T_4319_6;
  assign T_38374 = T_38373 & T_4319_5;
  assign T_38375 = T_38374 & T_4319_4;
  assign T_38376 = T_38375 & T_4319_3;
  assign T_38377 = T_38376 & T_4319_2;
  assign T_38378 = T_38377 & T_4319_1;
  assign T_38379 = T_38378 & T_4319_0;
  assign T_38390 = T_35573 & T_4324_21;
  assign T_38391 = T_38390 & T_4324_20;
  assign T_38392 = T_38391 & T_4324_19;
  assign T_38393 = T_38392 & T_4324_18;
  assign T_38394 = T_38393 & T_4324_17;
  assign T_38395 = T_38394 & T_4324_16;
  assign T_38396 = T_38395 & T_4324_15;
  assign T_38397 = T_38396 & T_4324_14;
  assign T_38398 = T_38397 & T_4324_13;
  assign T_38399 = T_38398 & T_4324_12;
  assign T_38400 = T_38399 & T_4324_11;
  assign T_38401 = T_38400 & T_4324_10;
  assign T_38402 = T_38401 & T_4324_9;
  assign T_38403 = T_38402 & T_4324_8;
  assign T_38404 = T_38403 & T_4324_7;
  assign T_38405 = T_38404 & T_4324_6;
  assign T_38406 = T_38405 & T_4324_5;
  assign T_38407 = T_38406 & T_4324_4;
  assign T_38408 = T_38407 & T_4324_3;
  assign T_38409 = T_38408 & T_4324_2;
  assign T_38410 = T_38409 & T_4324_1;
  assign T_38411 = T_38410 & T_4324_0;
  assign T_38422 = T_35605 & T_4329_21;
  assign T_38423 = T_38422 & T_4329_20;
  assign T_38424 = T_38423 & T_4329_19;
  assign T_38425 = T_38424 & T_4329_18;
  assign T_38426 = T_38425 & T_4329_17;
  assign T_38427 = T_38426 & T_4329_16;
  assign T_38428 = T_38427 & T_4329_15;
  assign T_38429 = T_38428 & T_4329_14;
  assign T_38430 = T_38429 & T_4329_13;
  assign T_38431 = T_38430 & T_4329_12;
  assign T_38432 = T_38431 & T_4329_11;
  assign T_38433 = T_38432 & T_4329_10;
  assign T_38434 = T_38433 & T_4329_9;
  assign T_38435 = T_38434 & T_4329_8;
  assign T_38436 = T_38435 & T_4329_7;
  assign T_38437 = T_38436 & T_4329_6;
  assign T_38438 = T_38437 & T_4329_5;
  assign T_38439 = T_38438 & T_4329_4;
  assign T_38440 = T_38439 & T_4329_3;
  assign T_38441 = T_38440 & T_4329_2;
  assign T_38442 = T_38441 & T_4329_1;
  assign T_38443 = T_38442 & T_4329_0;
  assign T_38454 = T_35637 & T_4334_21;
  assign T_38455 = T_38454 & T_4334_20;
  assign T_38456 = T_38455 & T_4334_19;
  assign T_38457 = T_38456 & T_4334_18;
  assign T_38458 = T_38457 & T_4334_17;
  assign T_38459 = T_38458 & T_4334_16;
  assign T_38460 = T_38459 & T_4334_15;
  assign T_38461 = T_38460 & T_4334_14;
  assign T_38462 = T_38461 & T_4334_13;
  assign T_38463 = T_38462 & T_4334_12;
  assign T_38464 = T_38463 & T_4334_11;
  assign T_38465 = T_38464 & T_4334_10;
  assign T_38466 = T_38465 & T_4334_9;
  assign T_38467 = T_38466 & T_4334_8;
  assign T_38468 = T_38467 & T_4334_7;
  assign T_38469 = T_38468 & T_4334_6;
  assign T_38470 = T_38469 & T_4334_5;
  assign T_38471 = T_38470 & T_4334_4;
  assign T_38472 = T_38471 & T_4334_3;
  assign T_38473 = T_38472 & T_4334_2;
  assign T_38474 = T_38473 & T_4334_1;
  assign T_38475 = T_38474 & T_4334_0;
  assign T_38485 = T_35540 & T_4319_22;
  assign T_38486 = T_38485 & T_4319_21;
  assign T_38487 = T_38486 & T_4319_20;
  assign T_38488 = T_38487 & T_4319_19;
  assign T_38489 = T_38488 & T_4319_18;
  assign T_38490 = T_38489 & T_4319_17;
  assign T_38491 = T_38490 & T_4319_16;
  assign T_38492 = T_38491 & T_4319_15;
  assign T_38493 = T_38492 & T_4319_14;
  assign T_38494 = T_38493 & T_4319_13;
  assign T_38495 = T_38494 & T_4319_12;
  assign T_38496 = T_38495 & T_4319_11;
  assign T_38497 = T_38496 & T_4319_10;
  assign T_38498 = T_38497 & T_4319_9;
  assign T_38499 = T_38498 & T_4319_8;
  assign T_38500 = T_38499 & T_4319_7;
  assign T_38501 = T_38500 & T_4319_6;
  assign T_38502 = T_38501 & T_4319_5;
  assign T_38503 = T_38502 & T_4319_4;
  assign T_38504 = T_38503 & T_4319_3;
  assign T_38505 = T_38504 & T_4319_2;
  assign T_38506 = T_38505 & T_4319_1;
  assign T_38507 = T_38506 & T_4319_0;
  assign T_38517 = T_35572 & T_4324_22;
  assign T_38518 = T_38517 & T_4324_21;
  assign T_38519 = T_38518 & T_4324_20;
  assign T_38520 = T_38519 & T_4324_19;
  assign T_38521 = T_38520 & T_4324_18;
  assign T_38522 = T_38521 & T_4324_17;
  assign T_38523 = T_38522 & T_4324_16;
  assign T_38524 = T_38523 & T_4324_15;
  assign T_38525 = T_38524 & T_4324_14;
  assign T_38526 = T_38525 & T_4324_13;
  assign T_38527 = T_38526 & T_4324_12;
  assign T_38528 = T_38527 & T_4324_11;
  assign T_38529 = T_38528 & T_4324_10;
  assign T_38530 = T_38529 & T_4324_9;
  assign T_38531 = T_38530 & T_4324_8;
  assign T_38532 = T_38531 & T_4324_7;
  assign T_38533 = T_38532 & T_4324_6;
  assign T_38534 = T_38533 & T_4324_5;
  assign T_38535 = T_38534 & T_4324_4;
  assign T_38536 = T_38535 & T_4324_3;
  assign T_38537 = T_38536 & T_4324_2;
  assign T_38538 = T_38537 & T_4324_1;
  assign T_38539 = T_38538 & T_4324_0;
  assign T_38549 = T_35604 & T_4329_22;
  assign T_38550 = T_38549 & T_4329_21;
  assign T_38551 = T_38550 & T_4329_20;
  assign T_38552 = T_38551 & T_4329_19;
  assign T_38553 = T_38552 & T_4329_18;
  assign T_38554 = T_38553 & T_4329_17;
  assign T_38555 = T_38554 & T_4329_16;
  assign T_38556 = T_38555 & T_4329_15;
  assign T_38557 = T_38556 & T_4329_14;
  assign T_38558 = T_38557 & T_4329_13;
  assign T_38559 = T_38558 & T_4329_12;
  assign T_38560 = T_38559 & T_4329_11;
  assign T_38561 = T_38560 & T_4329_10;
  assign T_38562 = T_38561 & T_4329_9;
  assign T_38563 = T_38562 & T_4329_8;
  assign T_38564 = T_38563 & T_4329_7;
  assign T_38565 = T_38564 & T_4329_6;
  assign T_38566 = T_38565 & T_4329_5;
  assign T_38567 = T_38566 & T_4329_4;
  assign T_38568 = T_38567 & T_4329_3;
  assign T_38569 = T_38568 & T_4329_2;
  assign T_38570 = T_38569 & T_4329_1;
  assign T_38571 = T_38570 & T_4329_0;
  assign T_38581 = T_35636 & T_4334_22;
  assign T_38582 = T_38581 & T_4334_21;
  assign T_38583 = T_38582 & T_4334_20;
  assign T_38584 = T_38583 & T_4334_19;
  assign T_38585 = T_38584 & T_4334_18;
  assign T_38586 = T_38585 & T_4334_17;
  assign T_38587 = T_38586 & T_4334_16;
  assign T_38588 = T_38587 & T_4334_15;
  assign T_38589 = T_38588 & T_4334_14;
  assign T_38590 = T_38589 & T_4334_13;
  assign T_38591 = T_38590 & T_4334_12;
  assign T_38592 = T_38591 & T_4334_11;
  assign T_38593 = T_38592 & T_4334_10;
  assign T_38594 = T_38593 & T_4334_9;
  assign T_38595 = T_38594 & T_4334_8;
  assign T_38596 = T_38595 & T_4334_7;
  assign T_38597 = T_38596 & T_4334_6;
  assign T_38598 = T_38597 & T_4334_5;
  assign T_38599 = T_38598 & T_4334_4;
  assign T_38600 = T_38599 & T_4334_3;
  assign T_38601 = T_38600 & T_4334_2;
  assign T_38602 = T_38601 & T_4334_1;
  assign T_38603 = T_38602 & T_4334_0;
  assign T_38612 = T_35539 & T_4319_23;
  assign T_38613 = T_38612 & T_4319_22;
  assign T_38614 = T_38613 & T_4319_21;
  assign T_38615 = T_38614 & T_4319_20;
  assign T_38616 = T_38615 & T_4319_19;
  assign T_38617 = T_38616 & T_4319_18;
  assign T_38618 = T_38617 & T_4319_17;
  assign T_38619 = T_38618 & T_4319_16;
  assign T_38620 = T_38619 & T_4319_15;
  assign T_38621 = T_38620 & T_4319_14;
  assign T_38622 = T_38621 & T_4319_13;
  assign T_38623 = T_38622 & T_4319_12;
  assign T_38624 = T_38623 & T_4319_11;
  assign T_38625 = T_38624 & T_4319_10;
  assign T_38626 = T_38625 & T_4319_9;
  assign T_38627 = T_38626 & T_4319_8;
  assign T_38628 = T_38627 & T_4319_7;
  assign T_38629 = T_38628 & T_4319_6;
  assign T_38630 = T_38629 & T_4319_5;
  assign T_38631 = T_38630 & T_4319_4;
  assign T_38632 = T_38631 & T_4319_3;
  assign T_38633 = T_38632 & T_4319_2;
  assign T_38634 = T_38633 & T_4319_1;
  assign T_38635 = T_38634 & T_4319_0;
  assign T_38644 = T_35571 & T_4324_23;
  assign T_38645 = T_38644 & T_4324_22;
  assign T_38646 = T_38645 & T_4324_21;
  assign T_38647 = T_38646 & T_4324_20;
  assign T_38648 = T_38647 & T_4324_19;
  assign T_38649 = T_38648 & T_4324_18;
  assign T_38650 = T_38649 & T_4324_17;
  assign T_38651 = T_38650 & T_4324_16;
  assign T_38652 = T_38651 & T_4324_15;
  assign T_38653 = T_38652 & T_4324_14;
  assign T_38654 = T_38653 & T_4324_13;
  assign T_38655 = T_38654 & T_4324_12;
  assign T_38656 = T_38655 & T_4324_11;
  assign T_38657 = T_38656 & T_4324_10;
  assign T_38658 = T_38657 & T_4324_9;
  assign T_38659 = T_38658 & T_4324_8;
  assign T_38660 = T_38659 & T_4324_7;
  assign T_38661 = T_38660 & T_4324_6;
  assign T_38662 = T_38661 & T_4324_5;
  assign T_38663 = T_38662 & T_4324_4;
  assign T_38664 = T_38663 & T_4324_3;
  assign T_38665 = T_38664 & T_4324_2;
  assign T_38666 = T_38665 & T_4324_1;
  assign T_38667 = T_38666 & T_4324_0;
  assign T_38676 = T_35603 & T_4329_23;
  assign T_38677 = T_38676 & T_4329_22;
  assign T_38678 = T_38677 & T_4329_21;
  assign T_38679 = T_38678 & T_4329_20;
  assign T_38680 = T_38679 & T_4329_19;
  assign T_38681 = T_38680 & T_4329_18;
  assign T_38682 = T_38681 & T_4329_17;
  assign T_38683 = T_38682 & T_4329_16;
  assign T_38684 = T_38683 & T_4329_15;
  assign T_38685 = T_38684 & T_4329_14;
  assign T_38686 = T_38685 & T_4329_13;
  assign T_38687 = T_38686 & T_4329_12;
  assign T_38688 = T_38687 & T_4329_11;
  assign T_38689 = T_38688 & T_4329_10;
  assign T_38690 = T_38689 & T_4329_9;
  assign T_38691 = T_38690 & T_4329_8;
  assign T_38692 = T_38691 & T_4329_7;
  assign T_38693 = T_38692 & T_4329_6;
  assign T_38694 = T_38693 & T_4329_5;
  assign T_38695 = T_38694 & T_4329_4;
  assign T_38696 = T_38695 & T_4329_3;
  assign T_38697 = T_38696 & T_4329_2;
  assign T_38698 = T_38697 & T_4329_1;
  assign T_38699 = T_38698 & T_4329_0;
  assign T_38708 = T_35635 & T_4334_23;
  assign T_38709 = T_38708 & T_4334_22;
  assign T_38710 = T_38709 & T_4334_21;
  assign T_38711 = T_38710 & T_4334_20;
  assign T_38712 = T_38711 & T_4334_19;
  assign T_38713 = T_38712 & T_4334_18;
  assign T_38714 = T_38713 & T_4334_17;
  assign T_38715 = T_38714 & T_4334_16;
  assign T_38716 = T_38715 & T_4334_15;
  assign T_38717 = T_38716 & T_4334_14;
  assign T_38718 = T_38717 & T_4334_13;
  assign T_38719 = T_38718 & T_4334_12;
  assign T_38720 = T_38719 & T_4334_11;
  assign T_38721 = T_38720 & T_4334_10;
  assign T_38722 = T_38721 & T_4334_9;
  assign T_38723 = T_38722 & T_4334_8;
  assign T_38724 = T_38723 & T_4334_7;
  assign T_38725 = T_38724 & T_4334_6;
  assign T_38726 = T_38725 & T_4334_5;
  assign T_38727 = T_38726 & T_4334_4;
  assign T_38728 = T_38727 & T_4334_3;
  assign T_38729 = T_38728 & T_4334_2;
  assign T_38730 = T_38729 & T_4334_1;
  assign T_38731 = T_38730 & T_4334_0;
  assign T_38739 = T_35538 & T_4319_24;
  assign T_38740 = T_38739 & T_4319_23;
  assign T_38741 = T_38740 & T_4319_22;
  assign T_38742 = T_38741 & T_4319_21;
  assign T_38743 = T_38742 & T_4319_20;
  assign T_38744 = T_38743 & T_4319_19;
  assign T_38745 = T_38744 & T_4319_18;
  assign T_38746 = T_38745 & T_4319_17;
  assign T_38747 = T_38746 & T_4319_16;
  assign T_38748 = T_38747 & T_4319_15;
  assign T_38749 = T_38748 & T_4319_14;
  assign T_38750 = T_38749 & T_4319_13;
  assign T_38751 = T_38750 & T_4319_12;
  assign T_38752 = T_38751 & T_4319_11;
  assign T_38753 = T_38752 & T_4319_10;
  assign T_38754 = T_38753 & T_4319_9;
  assign T_38755 = T_38754 & T_4319_8;
  assign T_38756 = T_38755 & T_4319_7;
  assign T_38757 = T_38756 & T_4319_6;
  assign T_38758 = T_38757 & T_4319_5;
  assign T_38759 = T_38758 & T_4319_4;
  assign T_38760 = T_38759 & T_4319_3;
  assign T_38761 = T_38760 & T_4319_2;
  assign T_38762 = T_38761 & T_4319_1;
  assign T_38763 = T_38762 & T_4319_0;
  assign T_38771 = T_35570 & T_4324_24;
  assign T_38772 = T_38771 & T_4324_23;
  assign T_38773 = T_38772 & T_4324_22;
  assign T_38774 = T_38773 & T_4324_21;
  assign T_38775 = T_38774 & T_4324_20;
  assign T_38776 = T_38775 & T_4324_19;
  assign T_38777 = T_38776 & T_4324_18;
  assign T_38778 = T_38777 & T_4324_17;
  assign T_38779 = T_38778 & T_4324_16;
  assign T_38780 = T_38779 & T_4324_15;
  assign T_38781 = T_38780 & T_4324_14;
  assign T_38782 = T_38781 & T_4324_13;
  assign T_38783 = T_38782 & T_4324_12;
  assign T_38784 = T_38783 & T_4324_11;
  assign T_38785 = T_38784 & T_4324_10;
  assign T_38786 = T_38785 & T_4324_9;
  assign T_38787 = T_38786 & T_4324_8;
  assign T_38788 = T_38787 & T_4324_7;
  assign T_38789 = T_38788 & T_4324_6;
  assign T_38790 = T_38789 & T_4324_5;
  assign T_38791 = T_38790 & T_4324_4;
  assign T_38792 = T_38791 & T_4324_3;
  assign T_38793 = T_38792 & T_4324_2;
  assign T_38794 = T_38793 & T_4324_1;
  assign T_38795 = T_38794 & T_4324_0;
  assign T_38803 = T_35602 & T_4329_24;
  assign T_38804 = T_38803 & T_4329_23;
  assign T_38805 = T_38804 & T_4329_22;
  assign T_38806 = T_38805 & T_4329_21;
  assign T_38807 = T_38806 & T_4329_20;
  assign T_38808 = T_38807 & T_4329_19;
  assign T_38809 = T_38808 & T_4329_18;
  assign T_38810 = T_38809 & T_4329_17;
  assign T_38811 = T_38810 & T_4329_16;
  assign T_38812 = T_38811 & T_4329_15;
  assign T_38813 = T_38812 & T_4329_14;
  assign T_38814 = T_38813 & T_4329_13;
  assign T_38815 = T_38814 & T_4329_12;
  assign T_38816 = T_38815 & T_4329_11;
  assign T_38817 = T_38816 & T_4329_10;
  assign T_38818 = T_38817 & T_4329_9;
  assign T_38819 = T_38818 & T_4329_8;
  assign T_38820 = T_38819 & T_4329_7;
  assign T_38821 = T_38820 & T_4329_6;
  assign T_38822 = T_38821 & T_4329_5;
  assign T_38823 = T_38822 & T_4329_4;
  assign T_38824 = T_38823 & T_4329_3;
  assign T_38825 = T_38824 & T_4329_2;
  assign T_38826 = T_38825 & T_4329_1;
  assign T_38827 = T_38826 & T_4329_0;
  assign T_38835 = T_35634 & T_4334_24;
  assign T_38836 = T_38835 & T_4334_23;
  assign T_38837 = T_38836 & T_4334_22;
  assign T_38838 = T_38837 & T_4334_21;
  assign T_38839 = T_38838 & T_4334_20;
  assign T_38840 = T_38839 & T_4334_19;
  assign T_38841 = T_38840 & T_4334_18;
  assign T_38842 = T_38841 & T_4334_17;
  assign T_38843 = T_38842 & T_4334_16;
  assign T_38844 = T_38843 & T_4334_15;
  assign T_38845 = T_38844 & T_4334_14;
  assign T_38846 = T_38845 & T_4334_13;
  assign T_38847 = T_38846 & T_4334_12;
  assign T_38848 = T_38847 & T_4334_11;
  assign T_38849 = T_38848 & T_4334_10;
  assign T_38850 = T_38849 & T_4334_9;
  assign T_38851 = T_38850 & T_4334_8;
  assign T_38852 = T_38851 & T_4334_7;
  assign T_38853 = T_38852 & T_4334_6;
  assign T_38854 = T_38853 & T_4334_5;
  assign T_38855 = T_38854 & T_4334_4;
  assign T_38856 = T_38855 & T_4334_3;
  assign T_38857 = T_38856 & T_4334_2;
  assign T_38858 = T_38857 & T_4334_1;
  assign T_38859 = T_38858 & T_4334_0;
  assign T_38866 = T_35537 & T_4319_25;
  assign T_38867 = T_38866 & T_4319_24;
  assign T_38868 = T_38867 & T_4319_23;
  assign T_38869 = T_38868 & T_4319_22;
  assign T_38870 = T_38869 & T_4319_21;
  assign T_38871 = T_38870 & T_4319_20;
  assign T_38872 = T_38871 & T_4319_19;
  assign T_38873 = T_38872 & T_4319_18;
  assign T_38874 = T_38873 & T_4319_17;
  assign T_38875 = T_38874 & T_4319_16;
  assign T_38876 = T_38875 & T_4319_15;
  assign T_38877 = T_38876 & T_4319_14;
  assign T_38878 = T_38877 & T_4319_13;
  assign T_38879 = T_38878 & T_4319_12;
  assign T_38880 = T_38879 & T_4319_11;
  assign T_38881 = T_38880 & T_4319_10;
  assign T_38882 = T_38881 & T_4319_9;
  assign T_38883 = T_38882 & T_4319_8;
  assign T_38884 = T_38883 & T_4319_7;
  assign T_38885 = T_38884 & T_4319_6;
  assign T_38886 = T_38885 & T_4319_5;
  assign T_38887 = T_38886 & T_4319_4;
  assign T_38888 = T_38887 & T_4319_3;
  assign T_38889 = T_38888 & T_4319_2;
  assign T_38890 = T_38889 & T_4319_1;
  assign T_38891 = T_38890 & T_4319_0;
  assign T_38898 = T_35569 & T_4324_25;
  assign T_38899 = T_38898 & T_4324_24;
  assign T_38900 = T_38899 & T_4324_23;
  assign T_38901 = T_38900 & T_4324_22;
  assign T_38902 = T_38901 & T_4324_21;
  assign T_38903 = T_38902 & T_4324_20;
  assign T_38904 = T_38903 & T_4324_19;
  assign T_38905 = T_38904 & T_4324_18;
  assign T_38906 = T_38905 & T_4324_17;
  assign T_38907 = T_38906 & T_4324_16;
  assign T_38908 = T_38907 & T_4324_15;
  assign T_38909 = T_38908 & T_4324_14;
  assign T_38910 = T_38909 & T_4324_13;
  assign T_38911 = T_38910 & T_4324_12;
  assign T_38912 = T_38911 & T_4324_11;
  assign T_38913 = T_38912 & T_4324_10;
  assign T_38914 = T_38913 & T_4324_9;
  assign T_38915 = T_38914 & T_4324_8;
  assign T_38916 = T_38915 & T_4324_7;
  assign T_38917 = T_38916 & T_4324_6;
  assign T_38918 = T_38917 & T_4324_5;
  assign T_38919 = T_38918 & T_4324_4;
  assign T_38920 = T_38919 & T_4324_3;
  assign T_38921 = T_38920 & T_4324_2;
  assign T_38922 = T_38921 & T_4324_1;
  assign T_38923 = T_38922 & T_4324_0;
  assign T_38930 = T_35601 & T_4329_25;
  assign T_38931 = T_38930 & T_4329_24;
  assign T_38932 = T_38931 & T_4329_23;
  assign T_38933 = T_38932 & T_4329_22;
  assign T_38934 = T_38933 & T_4329_21;
  assign T_38935 = T_38934 & T_4329_20;
  assign T_38936 = T_38935 & T_4329_19;
  assign T_38937 = T_38936 & T_4329_18;
  assign T_38938 = T_38937 & T_4329_17;
  assign T_38939 = T_38938 & T_4329_16;
  assign T_38940 = T_38939 & T_4329_15;
  assign T_38941 = T_38940 & T_4329_14;
  assign T_38942 = T_38941 & T_4329_13;
  assign T_38943 = T_38942 & T_4329_12;
  assign T_38944 = T_38943 & T_4329_11;
  assign T_38945 = T_38944 & T_4329_10;
  assign T_38946 = T_38945 & T_4329_9;
  assign T_38947 = T_38946 & T_4329_8;
  assign T_38948 = T_38947 & T_4329_7;
  assign T_38949 = T_38948 & T_4329_6;
  assign T_38950 = T_38949 & T_4329_5;
  assign T_38951 = T_38950 & T_4329_4;
  assign T_38952 = T_38951 & T_4329_3;
  assign T_38953 = T_38952 & T_4329_2;
  assign T_38954 = T_38953 & T_4329_1;
  assign T_38955 = T_38954 & T_4329_0;
  assign T_38962 = T_35633 & T_4334_25;
  assign T_38963 = T_38962 & T_4334_24;
  assign T_38964 = T_38963 & T_4334_23;
  assign T_38965 = T_38964 & T_4334_22;
  assign T_38966 = T_38965 & T_4334_21;
  assign T_38967 = T_38966 & T_4334_20;
  assign T_38968 = T_38967 & T_4334_19;
  assign T_38969 = T_38968 & T_4334_18;
  assign T_38970 = T_38969 & T_4334_17;
  assign T_38971 = T_38970 & T_4334_16;
  assign T_38972 = T_38971 & T_4334_15;
  assign T_38973 = T_38972 & T_4334_14;
  assign T_38974 = T_38973 & T_4334_13;
  assign T_38975 = T_38974 & T_4334_12;
  assign T_38976 = T_38975 & T_4334_11;
  assign T_38977 = T_38976 & T_4334_10;
  assign T_38978 = T_38977 & T_4334_9;
  assign T_38979 = T_38978 & T_4334_8;
  assign T_38980 = T_38979 & T_4334_7;
  assign T_38981 = T_38980 & T_4334_6;
  assign T_38982 = T_38981 & T_4334_5;
  assign T_38983 = T_38982 & T_4334_4;
  assign T_38984 = T_38983 & T_4334_3;
  assign T_38985 = T_38984 & T_4334_2;
  assign T_38986 = T_38985 & T_4334_1;
  assign T_38987 = T_38986 & T_4334_0;
  assign T_38993 = T_35536 & T_4319_26;
  assign T_38994 = T_38993 & T_4319_25;
  assign T_38995 = T_38994 & T_4319_24;
  assign T_38996 = T_38995 & T_4319_23;
  assign T_38997 = T_38996 & T_4319_22;
  assign T_38998 = T_38997 & T_4319_21;
  assign T_38999 = T_38998 & T_4319_20;
  assign T_39000 = T_38999 & T_4319_19;
  assign T_39001 = T_39000 & T_4319_18;
  assign T_39002 = T_39001 & T_4319_17;
  assign T_39003 = T_39002 & T_4319_16;
  assign T_39004 = T_39003 & T_4319_15;
  assign T_39005 = T_39004 & T_4319_14;
  assign T_39006 = T_39005 & T_4319_13;
  assign T_39007 = T_39006 & T_4319_12;
  assign T_39008 = T_39007 & T_4319_11;
  assign T_39009 = T_39008 & T_4319_10;
  assign T_39010 = T_39009 & T_4319_9;
  assign T_39011 = T_39010 & T_4319_8;
  assign T_39012 = T_39011 & T_4319_7;
  assign T_39013 = T_39012 & T_4319_6;
  assign T_39014 = T_39013 & T_4319_5;
  assign T_39015 = T_39014 & T_4319_4;
  assign T_39016 = T_39015 & T_4319_3;
  assign T_39017 = T_39016 & T_4319_2;
  assign T_39018 = T_39017 & T_4319_1;
  assign T_39019 = T_39018 & T_4319_0;
  assign T_39025 = T_35568 & T_4324_26;
  assign T_39026 = T_39025 & T_4324_25;
  assign T_39027 = T_39026 & T_4324_24;
  assign T_39028 = T_39027 & T_4324_23;
  assign T_39029 = T_39028 & T_4324_22;
  assign T_39030 = T_39029 & T_4324_21;
  assign T_39031 = T_39030 & T_4324_20;
  assign T_39032 = T_39031 & T_4324_19;
  assign T_39033 = T_39032 & T_4324_18;
  assign T_39034 = T_39033 & T_4324_17;
  assign T_39035 = T_39034 & T_4324_16;
  assign T_39036 = T_39035 & T_4324_15;
  assign T_39037 = T_39036 & T_4324_14;
  assign T_39038 = T_39037 & T_4324_13;
  assign T_39039 = T_39038 & T_4324_12;
  assign T_39040 = T_39039 & T_4324_11;
  assign T_39041 = T_39040 & T_4324_10;
  assign T_39042 = T_39041 & T_4324_9;
  assign T_39043 = T_39042 & T_4324_8;
  assign T_39044 = T_39043 & T_4324_7;
  assign T_39045 = T_39044 & T_4324_6;
  assign T_39046 = T_39045 & T_4324_5;
  assign T_39047 = T_39046 & T_4324_4;
  assign T_39048 = T_39047 & T_4324_3;
  assign T_39049 = T_39048 & T_4324_2;
  assign T_39050 = T_39049 & T_4324_1;
  assign T_39051 = T_39050 & T_4324_0;
  assign T_39057 = T_35600 & T_4329_26;
  assign T_39058 = T_39057 & T_4329_25;
  assign T_39059 = T_39058 & T_4329_24;
  assign T_39060 = T_39059 & T_4329_23;
  assign T_39061 = T_39060 & T_4329_22;
  assign T_39062 = T_39061 & T_4329_21;
  assign T_39063 = T_39062 & T_4329_20;
  assign T_39064 = T_39063 & T_4329_19;
  assign T_39065 = T_39064 & T_4329_18;
  assign T_39066 = T_39065 & T_4329_17;
  assign T_39067 = T_39066 & T_4329_16;
  assign T_39068 = T_39067 & T_4329_15;
  assign T_39069 = T_39068 & T_4329_14;
  assign T_39070 = T_39069 & T_4329_13;
  assign T_39071 = T_39070 & T_4329_12;
  assign T_39072 = T_39071 & T_4329_11;
  assign T_39073 = T_39072 & T_4329_10;
  assign T_39074 = T_39073 & T_4329_9;
  assign T_39075 = T_39074 & T_4329_8;
  assign T_39076 = T_39075 & T_4329_7;
  assign T_39077 = T_39076 & T_4329_6;
  assign T_39078 = T_39077 & T_4329_5;
  assign T_39079 = T_39078 & T_4329_4;
  assign T_39080 = T_39079 & T_4329_3;
  assign T_39081 = T_39080 & T_4329_2;
  assign T_39082 = T_39081 & T_4329_1;
  assign T_39083 = T_39082 & T_4329_0;
  assign T_39089 = T_35632 & T_4334_26;
  assign T_39090 = T_39089 & T_4334_25;
  assign T_39091 = T_39090 & T_4334_24;
  assign T_39092 = T_39091 & T_4334_23;
  assign T_39093 = T_39092 & T_4334_22;
  assign T_39094 = T_39093 & T_4334_21;
  assign T_39095 = T_39094 & T_4334_20;
  assign T_39096 = T_39095 & T_4334_19;
  assign T_39097 = T_39096 & T_4334_18;
  assign T_39098 = T_39097 & T_4334_17;
  assign T_39099 = T_39098 & T_4334_16;
  assign T_39100 = T_39099 & T_4334_15;
  assign T_39101 = T_39100 & T_4334_14;
  assign T_39102 = T_39101 & T_4334_13;
  assign T_39103 = T_39102 & T_4334_12;
  assign T_39104 = T_39103 & T_4334_11;
  assign T_39105 = T_39104 & T_4334_10;
  assign T_39106 = T_39105 & T_4334_9;
  assign T_39107 = T_39106 & T_4334_8;
  assign T_39108 = T_39107 & T_4334_7;
  assign T_39109 = T_39108 & T_4334_6;
  assign T_39110 = T_39109 & T_4334_5;
  assign T_39111 = T_39110 & T_4334_4;
  assign T_39112 = T_39111 & T_4334_3;
  assign T_39113 = T_39112 & T_4334_2;
  assign T_39114 = T_39113 & T_4334_1;
  assign T_39115 = T_39114 & T_4334_0;
  assign T_39120 = T_35535 & T_4319_27;
  assign T_39121 = T_39120 & T_4319_26;
  assign T_39122 = T_39121 & T_4319_25;
  assign T_39123 = T_39122 & T_4319_24;
  assign T_39124 = T_39123 & T_4319_23;
  assign T_39125 = T_39124 & T_4319_22;
  assign T_39126 = T_39125 & T_4319_21;
  assign T_39127 = T_39126 & T_4319_20;
  assign T_39128 = T_39127 & T_4319_19;
  assign T_39129 = T_39128 & T_4319_18;
  assign T_39130 = T_39129 & T_4319_17;
  assign T_39131 = T_39130 & T_4319_16;
  assign T_39132 = T_39131 & T_4319_15;
  assign T_39133 = T_39132 & T_4319_14;
  assign T_39134 = T_39133 & T_4319_13;
  assign T_39135 = T_39134 & T_4319_12;
  assign T_39136 = T_39135 & T_4319_11;
  assign T_39137 = T_39136 & T_4319_10;
  assign T_39138 = T_39137 & T_4319_9;
  assign T_39139 = T_39138 & T_4319_8;
  assign T_39140 = T_39139 & T_4319_7;
  assign T_39141 = T_39140 & T_4319_6;
  assign T_39142 = T_39141 & T_4319_5;
  assign T_39143 = T_39142 & T_4319_4;
  assign T_39144 = T_39143 & T_4319_3;
  assign T_39145 = T_39144 & T_4319_2;
  assign T_39146 = T_39145 & T_4319_1;
  assign T_39147 = T_39146 & T_4319_0;
  assign T_39152 = T_35567 & T_4324_27;
  assign T_39153 = T_39152 & T_4324_26;
  assign T_39154 = T_39153 & T_4324_25;
  assign T_39155 = T_39154 & T_4324_24;
  assign T_39156 = T_39155 & T_4324_23;
  assign T_39157 = T_39156 & T_4324_22;
  assign T_39158 = T_39157 & T_4324_21;
  assign T_39159 = T_39158 & T_4324_20;
  assign T_39160 = T_39159 & T_4324_19;
  assign T_39161 = T_39160 & T_4324_18;
  assign T_39162 = T_39161 & T_4324_17;
  assign T_39163 = T_39162 & T_4324_16;
  assign T_39164 = T_39163 & T_4324_15;
  assign T_39165 = T_39164 & T_4324_14;
  assign T_39166 = T_39165 & T_4324_13;
  assign T_39167 = T_39166 & T_4324_12;
  assign T_39168 = T_39167 & T_4324_11;
  assign T_39169 = T_39168 & T_4324_10;
  assign T_39170 = T_39169 & T_4324_9;
  assign T_39171 = T_39170 & T_4324_8;
  assign T_39172 = T_39171 & T_4324_7;
  assign T_39173 = T_39172 & T_4324_6;
  assign T_39174 = T_39173 & T_4324_5;
  assign T_39175 = T_39174 & T_4324_4;
  assign T_39176 = T_39175 & T_4324_3;
  assign T_39177 = T_39176 & T_4324_2;
  assign T_39178 = T_39177 & T_4324_1;
  assign T_39179 = T_39178 & T_4324_0;
  assign T_39184 = T_35599 & T_4329_27;
  assign T_39185 = T_39184 & T_4329_26;
  assign T_39186 = T_39185 & T_4329_25;
  assign T_39187 = T_39186 & T_4329_24;
  assign T_39188 = T_39187 & T_4329_23;
  assign T_39189 = T_39188 & T_4329_22;
  assign T_39190 = T_39189 & T_4329_21;
  assign T_39191 = T_39190 & T_4329_20;
  assign T_39192 = T_39191 & T_4329_19;
  assign T_39193 = T_39192 & T_4329_18;
  assign T_39194 = T_39193 & T_4329_17;
  assign T_39195 = T_39194 & T_4329_16;
  assign T_39196 = T_39195 & T_4329_15;
  assign T_39197 = T_39196 & T_4329_14;
  assign T_39198 = T_39197 & T_4329_13;
  assign T_39199 = T_39198 & T_4329_12;
  assign T_39200 = T_39199 & T_4329_11;
  assign T_39201 = T_39200 & T_4329_10;
  assign T_39202 = T_39201 & T_4329_9;
  assign T_39203 = T_39202 & T_4329_8;
  assign T_39204 = T_39203 & T_4329_7;
  assign T_39205 = T_39204 & T_4329_6;
  assign T_39206 = T_39205 & T_4329_5;
  assign T_39207 = T_39206 & T_4329_4;
  assign T_39208 = T_39207 & T_4329_3;
  assign T_39209 = T_39208 & T_4329_2;
  assign T_39210 = T_39209 & T_4329_1;
  assign T_39211 = T_39210 & T_4329_0;
  assign T_39216 = T_35631 & T_4334_27;
  assign T_39217 = T_39216 & T_4334_26;
  assign T_39218 = T_39217 & T_4334_25;
  assign T_39219 = T_39218 & T_4334_24;
  assign T_39220 = T_39219 & T_4334_23;
  assign T_39221 = T_39220 & T_4334_22;
  assign T_39222 = T_39221 & T_4334_21;
  assign T_39223 = T_39222 & T_4334_20;
  assign T_39224 = T_39223 & T_4334_19;
  assign T_39225 = T_39224 & T_4334_18;
  assign T_39226 = T_39225 & T_4334_17;
  assign T_39227 = T_39226 & T_4334_16;
  assign T_39228 = T_39227 & T_4334_15;
  assign T_39229 = T_39228 & T_4334_14;
  assign T_39230 = T_39229 & T_4334_13;
  assign T_39231 = T_39230 & T_4334_12;
  assign T_39232 = T_39231 & T_4334_11;
  assign T_39233 = T_39232 & T_4334_10;
  assign T_39234 = T_39233 & T_4334_9;
  assign T_39235 = T_39234 & T_4334_8;
  assign T_39236 = T_39235 & T_4334_7;
  assign T_39237 = T_39236 & T_4334_6;
  assign T_39238 = T_39237 & T_4334_5;
  assign T_39239 = T_39238 & T_4334_4;
  assign T_39240 = T_39239 & T_4334_3;
  assign T_39241 = T_39240 & T_4334_2;
  assign T_39242 = T_39241 & T_4334_1;
  assign T_39243 = T_39242 & T_4334_0;
  assign T_39247 = T_35534 & T_4319_28;
  assign T_39248 = T_39247 & T_4319_27;
  assign T_39249 = T_39248 & T_4319_26;
  assign T_39250 = T_39249 & T_4319_25;
  assign T_39251 = T_39250 & T_4319_24;
  assign T_39252 = T_39251 & T_4319_23;
  assign T_39253 = T_39252 & T_4319_22;
  assign T_39254 = T_39253 & T_4319_21;
  assign T_39255 = T_39254 & T_4319_20;
  assign T_39256 = T_39255 & T_4319_19;
  assign T_39257 = T_39256 & T_4319_18;
  assign T_39258 = T_39257 & T_4319_17;
  assign T_39259 = T_39258 & T_4319_16;
  assign T_39260 = T_39259 & T_4319_15;
  assign T_39261 = T_39260 & T_4319_14;
  assign T_39262 = T_39261 & T_4319_13;
  assign T_39263 = T_39262 & T_4319_12;
  assign T_39264 = T_39263 & T_4319_11;
  assign T_39265 = T_39264 & T_4319_10;
  assign T_39266 = T_39265 & T_4319_9;
  assign T_39267 = T_39266 & T_4319_8;
  assign T_39268 = T_39267 & T_4319_7;
  assign T_39269 = T_39268 & T_4319_6;
  assign T_39270 = T_39269 & T_4319_5;
  assign T_39271 = T_39270 & T_4319_4;
  assign T_39272 = T_39271 & T_4319_3;
  assign T_39273 = T_39272 & T_4319_2;
  assign T_39274 = T_39273 & T_4319_1;
  assign T_39275 = T_39274 & T_4319_0;
  assign T_39279 = T_35566 & T_4324_28;
  assign T_39280 = T_39279 & T_4324_27;
  assign T_39281 = T_39280 & T_4324_26;
  assign T_39282 = T_39281 & T_4324_25;
  assign T_39283 = T_39282 & T_4324_24;
  assign T_39284 = T_39283 & T_4324_23;
  assign T_39285 = T_39284 & T_4324_22;
  assign T_39286 = T_39285 & T_4324_21;
  assign T_39287 = T_39286 & T_4324_20;
  assign T_39288 = T_39287 & T_4324_19;
  assign T_39289 = T_39288 & T_4324_18;
  assign T_39290 = T_39289 & T_4324_17;
  assign T_39291 = T_39290 & T_4324_16;
  assign T_39292 = T_39291 & T_4324_15;
  assign T_39293 = T_39292 & T_4324_14;
  assign T_39294 = T_39293 & T_4324_13;
  assign T_39295 = T_39294 & T_4324_12;
  assign T_39296 = T_39295 & T_4324_11;
  assign T_39297 = T_39296 & T_4324_10;
  assign T_39298 = T_39297 & T_4324_9;
  assign T_39299 = T_39298 & T_4324_8;
  assign T_39300 = T_39299 & T_4324_7;
  assign T_39301 = T_39300 & T_4324_6;
  assign T_39302 = T_39301 & T_4324_5;
  assign T_39303 = T_39302 & T_4324_4;
  assign T_39304 = T_39303 & T_4324_3;
  assign T_39305 = T_39304 & T_4324_2;
  assign T_39306 = T_39305 & T_4324_1;
  assign T_39307 = T_39306 & T_4324_0;
  assign T_39311 = T_35598 & T_4329_28;
  assign T_39312 = T_39311 & T_4329_27;
  assign T_39313 = T_39312 & T_4329_26;
  assign T_39314 = T_39313 & T_4329_25;
  assign T_39315 = T_39314 & T_4329_24;
  assign T_39316 = T_39315 & T_4329_23;
  assign T_39317 = T_39316 & T_4329_22;
  assign T_39318 = T_39317 & T_4329_21;
  assign T_39319 = T_39318 & T_4329_20;
  assign T_39320 = T_39319 & T_4329_19;
  assign T_39321 = T_39320 & T_4329_18;
  assign T_39322 = T_39321 & T_4329_17;
  assign T_39323 = T_39322 & T_4329_16;
  assign T_39324 = T_39323 & T_4329_15;
  assign T_39325 = T_39324 & T_4329_14;
  assign T_39326 = T_39325 & T_4329_13;
  assign T_39327 = T_39326 & T_4329_12;
  assign T_39328 = T_39327 & T_4329_11;
  assign T_39329 = T_39328 & T_4329_10;
  assign T_39330 = T_39329 & T_4329_9;
  assign T_39331 = T_39330 & T_4329_8;
  assign T_39332 = T_39331 & T_4329_7;
  assign T_39333 = T_39332 & T_4329_6;
  assign T_39334 = T_39333 & T_4329_5;
  assign T_39335 = T_39334 & T_4329_4;
  assign T_39336 = T_39335 & T_4329_3;
  assign T_39337 = T_39336 & T_4329_2;
  assign T_39338 = T_39337 & T_4329_1;
  assign T_39339 = T_39338 & T_4329_0;
  assign T_39343 = T_35630 & T_4334_28;
  assign T_39344 = T_39343 & T_4334_27;
  assign T_39345 = T_39344 & T_4334_26;
  assign T_39346 = T_39345 & T_4334_25;
  assign T_39347 = T_39346 & T_4334_24;
  assign T_39348 = T_39347 & T_4334_23;
  assign T_39349 = T_39348 & T_4334_22;
  assign T_39350 = T_39349 & T_4334_21;
  assign T_39351 = T_39350 & T_4334_20;
  assign T_39352 = T_39351 & T_4334_19;
  assign T_39353 = T_39352 & T_4334_18;
  assign T_39354 = T_39353 & T_4334_17;
  assign T_39355 = T_39354 & T_4334_16;
  assign T_39356 = T_39355 & T_4334_15;
  assign T_39357 = T_39356 & T_4334_14;
  assign T_39358 = T_39357 & T_4334_13;
  assign T_39359 = T_39358 & T_4334_12;
  assign T_39360 = T_39359 & T_4334_11;
  assign T_39361 = T_39360 & T_4334_10;
  assign T_39362 = T_39361 & T_4334_9;
  assign T_39363 = T_39362 & T_4334_8;
  assign T_39364 = T_39363 & T_4334_7;
  assign T_39365 = T_39364 & T_4334_6;
  assign T_39366 = T_39365 & T_4334_5;
  assign T_39367 = T_39366 & T_4334_4;
  assign T_39368 = T_39367 & T_4334_3;
  assign T_39369 = T_39368 & T_4334_2;
  assign T_39370 = T_39369 & T_4334_1;
  assign T_39371 = T_39370 & T_4334_0;
  assign T_39374 = T_35533 & T_4319_29;
  assign T_39375 = T_39374 & T_4319_28;
  assign T_39376 = T_39375 & T_4319_27;
  assign T_39377 = T_39376 & T_4319_26;
  assign T_39378 = T_39377 & T_4319_25;
  assign T_39379 = T_39378 & T_4319_24;
  assign T_39380 = T_39379 & T_4319_23;
  assign T_39381 = T_39380 & T_4319_22;
  assign T_39382 = T_39381 & T_4319_21;
  assign T_39383 = T_39382 & T_4319_20;
  assign T_39384 = T_39383 & T_4319_19;
  assign T_39385 = T_39384 & T_4319_18;
  assign T_39386 = T_39385 & T_4319_17;
  assign T_39387 = T_39386 & T_4319_16;
  assign T_39388 = T_39387 & T_4319_15;
  assign T_39389 = T_39388 & T_4319_14;
  assign T_39390 = T_39389 & T_4319_13;
  assign T_39391 = T_39390 & T_4319_12;
  assign T_39392 = T_39391 & T_4319_11;
  assign T_39393 = T_39392 & T_4319_10;
  assign T_39394 = T_39393 & T_4319_9;
  assign T_39395 = T_39394 & T_4319_8;
  assign T_39396 = T_39395 & T_4319_7;
  assign T_39397 = T_39396 & T_4319_6;
  assign T_39398 = T_39397 & T_4319_5;
  assign T_39399 = T_39398 & T_4319_4;
  assign T_39400 = T_39399 & T_4319_3;
  assign T_39401 = T_39400 & T_4319_2;
  assign T_39402 = T_39401 & T_4319_1;
  assign T_39403 = T_39402 & T_4319_0;
  assign T_39406 = T_35565 & T_4324_29;
  assign T_39407 = T_39406 & T_4324_28;
  assign T_39408 = T_39407 & T_4324_27;
  assign T_39409 = T_39408 & T_4324_26;
  assign T_39410 = T_39409 & T_4324_25;
  assign T_39411 = T_39410 & T_4324_24;
  assign T_39412 = T_39411 & T_4324_23;
  assign T_39413 = T_39412 & T_4324_22;
  assign T_39414 = T_39413 & T_4324_21;
  assign T_39415 = T_39414 & T_4324_20;
  assign T_39416 = T_39415 & T_4324_19;
  assign T_39417 = T_39416 & T_4324_18;
  assign T_39418 = T_39417 & T_4324_17;
  assign T_39419 = T_39418 & T_4324_16;
  assign T_39420 = T_39419 & T_4324_15;
  assign T_39421 = T_39420 & T_4324_14;
  assign T_39422 = T_39421 & T_4324_13;
  assign T_39423 = T_39422 & T_4324_12;
  assign T_39424 = T_39423 & T_4324_11;
  assign T_39425 = T_39424 & T_4324_10;
  assign T_39426 = T_39425 & T_4324_9;
  assign T_39427 = T_39426 & T_4324_8;
  assign T_39428 = T_39427 & T_4324_7;
  assign T_39429 = T_39428 & T_4324_6;
  assign T_39430 = T_39429 & T_4324_5;
  assign T_39431 = T_39430 & T_4324_4;
  assign T_39432 = T_39431 & T_4324_3;
  assign T_39433 = T_39432 & T_4324_2;
  assign T_39434 = T_39433 & T_4324_1;
  assign T_39435 = T_39434 & T_4324_0;
  assign T_39438 = T_35597 & T_4329_29;
  assign T_39439 = T_39438 & T_4329_28;
  assign T_39440 = T_39439 & T_4329_27;
  assign T_39441 = T_39440 & T_4329_26;
  assign T_39442 = T_39441 & T_4329_25;
  assign T_39443 = T_39442 & T_4329_24;
  assign T_39444 = T_39443 & T_4329_23;
  assign T_39445 = T_39444 & T_4329_22;
  assign T_39446 = T_39445 & T_4329_21;
  assign T_39447 = T_39446 & T_4329_20;
  assign T_39448 = T_39447 & T_4329_19;
  assign T_39449 = T_39448 & T_4329_18;
  assign T_39450 = T_39449 & T_4329_17;
  assign T_39451 = T_39450 & T_4329_16;
  assign T_39452 = T_39451 & T_4329_15;
  assign T_39453 = T_39452 & T_4329_14;
  assign T_39454 = T_39453 & T_4329_13;
  assign T_39455 = T_39454 & T_4329_12;
  assign T_39456 = T_39455 & T_4329_11;
  assign T_39457 = T_39456 & T_4329_10;
  assign T_39458 = T_39457 & T_4329_9;
  assign T_39459 = T_39458 & T_4329_8;
  assign T_39460 = T_39459 & T_4329_7;
  assign T_39461 = T_39460 & T_4329_6;
  assign T_39462 = T_39461 & T_4329_5;
  assign T_39463 = T_39462 & T_4329_4;
  assign T_39464 = T_39463 & T_4329_3;
  assign T_39465 = T_39464 & T_4329_2;
  assign T_39466 = T_39465 & T_4329_1;
  assign T_39467 = T_39466 & T_4329_0;
  assign T_39470 = T_35629 & T_4334_29;
  assign T_39471 = T_39470 & T_4334_28;
  assign T_39472 = T_39471 & T_4334_27;
  assign T_39473 = T_39472 & T_4334_26;
  assign T_39474 = T_39473 & T_4334_25;
  assign T_39475 = T_39474 & T_4334_24;
  assign T_39476 = T_39475 & T_4334_23;
  assign T_39477 = T_39476 & T_4334_22;
  assign T_39478 = T_39477 & T_4334_21;
  assign T_39479 = T_39478 & T_4334_20;
  assign T_39480 = T_39479 & T_4334_19;
  assign T_39481 = T_39480 & T_4334_18;
  assign T_39482 = T_39481 & T_4334_17;
  assign T_39483 = T_39482 & T_4334_16;
  assign T_39484 = T_39483 & T_4334_15;
  assign T_39485 = T_39484 & T_4334_14;
  assign T_39486 = T_39485 & T_4334_13;
  assign T_39487 = T_39486 & T_4334_12;
  assign T_39488 = T_39487 & T_4334_11;
  assign T_39489 = T_39488 & T_4334_10;
  assign T_39490 = T_39489 & T_4334_9;
  assign T_39491 = T_39490 & T_4334_8;
  assign T_39492 = T_39491 & T_4334_7;
  assign T_39493 = T_39492 & T_4334_6;
  assign T_39494 = T_39493 & T_4334_5;
  assign T_39495 = T_39494 & T_4334_4;
  assign T_39496 = T_39495 & T_4334_3;
  assign T_39497 = T_39496 & T_4334_2;
  assign T_39498 = T_39497 & T_4334_1;
  assign T_39499 = T_39498 & T_4334_0;
  assign T_39501 = T_26576 & T_4319_30;
  assign T_39502 = T_39501 & T_4319_29;
  assign T_39503 = T_39502 & T_4319_28;
  assign T_39504 = T_39503 & T_4319_27;
  assign T_39505 = T_39504 & T_4319_26;
  assign T_39506 = T_39505 & T_4319_25;
  assign T_39507 = T_39506 & T_4319_24;
  assign T_39508 = T_39507 & T_4319_23;
  assign T_39509 = T_39508 & T_4319_22;
  assign T_39510 = T_39509 & T_4319_21;
  assign T_39511 = T_39510 & T_4319_20;
  assign T_39512 = T_39511 & T_4319_19;
  assign T_39513 = T_39512 & T_4319_18;
  assign T_39514 = T_39513 & T_4319_17;
  assign T_39515 = T_39514 & T_4319_16;
  assign T_39516 = T_39515 & T_4319_15;
  assign T_39517 = T_39516 & T_4319_14;
  assign T_39518 = T_39517 & T_4319_13;
  assign T_39519 = T_39518 & T_4319_12;
  assign T_39520 = T_39519 & T_4319_11;
  assign T_39521 = T_39520 & T_4319_10;
  assign T_39522 = T_39521 & T_4319_9;
  assign T_39523 = T_39522 & T_4319_8;
  assign T_39524 = T_39523 & T_4319_7;
  assign T_39525 = T_39524 & T_4319_6;
  assign T_39526 = T_39525 & T_4319_5;
  assign T_39527 = T_39526 & T_4319_4;
  assign T_39528 = T_39527 & T_4319_3;
  assign T_39529 = T_39528 & T_4319_2;
  assign T_39530 = T_39529 & T_4319_1;
  assign T_39531 = T_39530 & T_4319_0;
  assign T_39533 = T_26582 & T_4324_30;
  assign T_39534 = T_39533 & T_4324_29;
  assign T_39535 = T_39534 & T_4324_28;
  assign T_39536 = T_39535 & T_4324_27;
  assign T_39537 = T_39536 & T_4324_26;
  assign T_39538 = T_39537 & T_4324_25;
  assign T_39539 = T_39538 & T_4324_24;
  assign T_39540 = T_39539 & T_4324_23;
  assign T_39541 = T_39540 & T_4324_22;
  assign T_39542 = T_39541 & T_4324_21;
  assign T_39543 = T_39542 & T_4324_20;
  assign T_39544 = T_39543 & T_4324_19;
  assign T_39545 = T_39544 & T_4324_18;
  assign T_39546 = T_39545 & T_4324_17;
  assign T_39547 = T_39546 & T_4324_16;
  assign T_39548 = T_39547 & T_4324_15;
  assign T_39549 = T_39548 & T_4324_14;
  assign T_39550 = T_39549 & T_4324_13;
  assign T_39551 = T_39550 & T_4324_12;
  assign T_39552 = T_39551 & T_4324_11;
  assign T_39553 = T_39552 & T_4324_10;
  assign T_39554 = T_39553 & T_4324_9;
  assign T_39555 = T_39554 & T_4324_8;
  assign T_39556 = T_39555 & T_4324_7;
  assign T_39557 = T_39556 & T_4324_6;
  assign T_39558 = T_39557 & T_4324_5;
  assign T_39559 = T_39558 & T_4324_4;
  assign T_39560 = T_39559 & T_4324_3;
  assign T_39561 = T_39560 & T_4324_2;
  assign T_39562 = T_39561 & T_4324_1;
  assign T_39563 = T_39562 & T_4324_0;
  assign T_39565 = T_26586 & T_4329_30;
  assign T_39566 = T_39565 & T_4329_29;
  assign T_39567 = T_39566 & T_4329_28;
  assign T_39568 = T_39567 & T_4329_27;
  assign T_39569 = T_39568 & T_4329_26;
  assign T_39570 = T_39569 & T_4329_25;
  assign T_39571 = T_39570 & T_4329_24;
  assign T_39572 = T_39571 & T_4329_23;
  assign T_39573 = T_39572 & T_4329_22;
  assign T_39574 = T_39573 & T_4329_21;
  assign T_39575 = T_39574 & T_4329_20;
  assign T_39576 = T_39575 & T_4329_19;
  assign T_39577 = T_39576 & T_4329_18;
  assign T_39578 = T_39577 & T_4329_17;
  assign T_39579 = T_39578 & T_4329_16;
  assign T_39580 = T_39579 & T_4329_15;
  assign T_39581 = T_39580 & T_4329_14;
  assign T_39582 = T_39581 & T_4329_13;
  assign T_39583 = T_39582 & T_4329_12;
  assign T_39584 = T_39583 & T_4329_11;
  assign T_39585 = T_39584 & T_4329_10;
  assign T_39586 = T_39585 & T_4329_9;
  assign T_39587 = T_39586 & T_4329_8;
  assign T_39588 = T_39587 & T_4329_7;
  assign T_39589 = T_39588 & T_4329_6;
  assign T_39590 = T_39589 & T_4329_5;
  assign T_39591 = T_39590 & T_4329_4;
  assign T_39592 = T_39591 & T_4329_3;
  assign T_39593 = T_39592 & T_4329_2;
  assign T_39594 = T_39593 & T_4329_1;
  assign T_39595 = T_39594 & T_4329_0;
  assign T_39597 = T_26592 & T_4334_30;
  assign T_39598 = T_39597 & T_4334_29;
  assign T_39599 = T_39598 & T_4334_28;
  assign T_39600 = T_39599 & T_4334_27;
  assign T_39601 = T_39600 & T_4334_26;
  assign T_39602 = T_39601 & T_4334_25;
  assign T_39603 = T_39602 & T_4334_24;
  assign T_39604 = T_39603 & T_4334_23;
  assign T_39605 = T_39604 & T_4334_22;
  assign T_39606 = T_39605 & T_4334_21;
  assign T_39607 = T_39606 & T_4334_20;
  assign T_39608 = T_39607 & T_4334_19;
  assign T_39609 = T_39608 & T_4334_18;
  assign T_39610 = T_39609 & T_4334_17;
  assign T_39611 = T_39610 & T_4334_16;
  assign T_39612 = T_39611 & T_4334_15;
  assign T_39613 = T_39612 & T_4334_14;
  assign T_39614 = T_39613 & T_4334_13;
  assign T_39615 = T_39614 & T_4334_12;
  assign T_39616 = T_39615 & T_4334_11;
  assign T_39617 = T_39616 & T_4334_10;
  assign T_39618 = T_39617 & T_4334_9;
  assign T_39619 = T_39618 & T_4334_8;
  assign T_39620 = T_39619 & T_4334_7;
  assign T_39621 = T_39620 & T_4334_6;
  assign T_39622 = T_39621 & T_4334_5;
  assign T_39623 = T_39622 & T_4334_4;
  assign T_39624 = T_39623 & T_4334_3;
  assign T_39625 = T_39624 & T_4334_2;
  assign T_39626 = T_39625 & T_4334_1;
  assign T_39627 = T_39626 & T_4334_0;
  assign T_39665 = T_27876 & T_4319_60;
  assign T_39666 = T_39665 & T_4319_59;
  assign T_39667 = T_39666 & T_4319_58;
  assign T_39668 = T_39667 & T_4319_57;
  assign T_39669 = T_39668 & T_4319_56;
  assign T_39670 = T_39669 & T_4319_55;
  assign T_39671 = T_39670 & T_4319_54;
  assign T_39672 = T_39671 & T_4319_53;
  assign T_39673 = T_39672 & T_4319_52;
  assign T_39674 = T_39673 & T_4319_51;
  assign T_39675 = T_39674 & T_4319_50;
  assign T_39676 = T_39675 & T_4319_49;
  assign T_39677 = T_39676 & T_4319_48;
  assign T_39678 = T_39677 & T_4319_47;
  assign T_39679 = T_39678 & T_4319_46;
  assign T_39680 = T_39679 & T_4319_45;
  assign T_39681 = T_39680 & T_4319_44;
  assign T_39682 = T_39681 & T_4319_43;
  assign T_39683 = T_39682 & T_4319_42;
  assign T_39685 = T_27882 & T_4324_60;
  assign T_39686 = T_39685 & T_4324_59;
  assign T_39687 = T_39686 & T_4324_58;
  assign T_39688 = T_39687 & T_4324_57;
  assign T_39689 = T_39688 & T_4324_56;
  assign T_39690 = T_39689 & T_4324_55;
  assign T_39691 = T_39690 & T_4324_54;
  assign T_39692 = T_39691 & T_4324_53;
  assign T_39693 = T_39692 & T_4324_52;
  assign T_39694 = T_39693 & T_4324_51;
  assign T_39695 = T_39694 & T_4324_50;
  assign T_39696 = T_39695 & T_4324_49;
  assign T_39697 = T_39696 & T_4324_48;
  assign T_39698 = T_39697 & T_4324_47;
  assign T_39699 = T_39698 & T_4324_46;
  assign T_39700 = T_39699 & T_4324_45;
  assign T_39701 = T_39700 & T_4324_44;
  assign T_39702 = T_39701 & T_4324_43;
  assign T_39703 = T_39702 & T_4324_42;
  assign T_39705 = T_27886 & T_4329_60;
  assign T_39706 = T_39705 & T_4329_59;
  assign T_39707 = T_39706 & T_4329_58;
  assign T_39708 = T_39707 & T_4329_57;
  assign T_39709 = T_39708 & T_4329_56;
  assign T_39710 = T_39709 & T_4329_55;
  assign T_39711 = T_39710 & T_4329_54;
  assign T_39712 = T_39711 & T_4329_53;
  assign T_39713 = T_39712 & T_4329_52;
  assign T_39714 = T_39713 & T_4329_51;
  assign T_39715 = T_39714 & T_4329_50;
  assign T_39716 = T_39715 & T_4329_49;
  assign T_39717 = T_39716 & T_4329_48;
  assign T_39718 = T_39717 & T_4329_47;
  assign T_39719 = T_39718 & T_4329_46;
  assign T_39720 = T_39719 & T_4329_45;
  assign T_39721 = T_39720 & T_4329_44;
  assign T_39722 = T_39721 & T_4329_43;
  assign T_39723 = T_39722 & T_4329_42;
  assign T_39725 = T_27892 & T_4334_60;
  assign T_39726 = T_39725 & T_4334_59;
  assign T_39727 = T_39726 & T_4334_58;
  assign T_39728 = T_39727 & T_4334_57;
  assign T_39729 = T_39728 & T_4334_56;
  assign T_39730 = T_39729 & T_4334_55;
  assign T_39731 = T_39730 & T_4334_54;
  assign T_39732 = T_39731 & T_4334_53;
  assign T_39733 = T_39732 & T_4334_52;
  assign T_39734 = T_39733 & T_4334_51;
  assign T_39735 = T_39734 & T_4334_50;
  assign T_39736 = T_39735 & T_4334_49;
  assign T_39737 = T_39736 & T_4334_48;
  assign T_39738 = T_39737 & T_4334_47;
  assign T_39739 = T_39738 & T_4334_46;
  assign T_39740 = T_39739 & T_4334_45;
  assign T_39741 = T_39740 & T_4334_44;
  assign T_39742 = T_39741 & T_4334_43;
  assign T_39743 = T_39742 & T_4334_42;
  assign T_39763 = T_39682 & T_4319_41;
  assign T_39783 = T_39702 & T_4324_41;
  assign T_39803 = T_39722 & T_4329_41;
  assign T_39823 = T_39742 & T_4334_41;
  assign T_39842 = T_39681 & T_4319_42;
  assign T_39843 = T_39842 & T_4319_41;
  assign T_39862 = T_39701 & T_4324_42;
  assign T_39863 = T_39862 & T_4324_41;
  assign T_39882 = T_39721 & T_4329_42;
  assign T_39883 = T_39882 & T_4329_41;
  assign T_39902 = T_39741 & T_4334_42;
  assign T_39903 = T_39902 & T_4334_41;
  assign T_39921 = T_39680 & T_4319_43;
  assign T_39922 = T_39921 & T_4319_42;
  assign T_39923 = T_39922 & T_4319_41;
  assign T_39941 = T_39700 & T_4324_43;
  assign T_39942 = T_39941 & T_4324_42;
  assign T_39943 = T_39942 & T_4324_41;
  assign T_39961 = T_39720 & T_4329_43;
  assign T_39962 = T_39961 & T_4329_42;
  assign T_39963 = T_39962 & T_4329_41;
  assign T_39981 = T_39740 & T_4334_43;
  assign T_39982 = T_39981 & T_4334_42;
  assign T_39983 = T_39982 & T_4334_41;
  assign T_40000 = T_39679 & T_4319_44;
  assign T_40001 = T_40000 & T_4319_43;
  assign T_40002 = T_40001 & T_4319_42;
  assign T_40003 = T_40002 & T_4319_41;
  assign T_40020 = T_39699 & T_4324_44;
  assign T_40021 = T_40020 & T_4324_43;
  assign T_40022 = T_40021 & T_4324_42;
  assign T_40023 = T_40022 & T_4324_41;
  assign T_40040 = T_39719 & T_4329_44;
  assign T_40041 = T_40040 & T_4329_43;
  assign T_40042 = T_40041 & T_4329_42;
  assign T_40043 = T_40042 & T_4329_41;
  assign T_40060 = T_39739 & T_4334_44;
  assign T_40061 = T_40060 & T_4334_43;
  assign T_40062 = T_40061 & T_4334_42;
  assign T_40063 = T_40062 & T_4334_41;
  assign T_40079 = T_39678 & T_4319_45;
  assign T_40080 = T_40079 & T_4319_44;
  assign T_40081 = T_40080 & T_4319_43;
  assign T_40082 = T_40081 & T_4319_42;
  assign T_40083 = T_40082 & T_4319_41;
  assign T_40099 = T_39698 & T_4324_45;
  assign T_40100 = T_40099 & T_4324_44;
  assign T_40101 = T_40100 & T_4324_43;
  assign T_40102 = T_40101 & T_4324_42;
  assign T_40103 = T_40102 & T_4324_41;
  assign T_40119 = T_39718 & T_4329_45;
  assign T_40120 = T_40119 & T_4329_44;
  assign T_40121 = T_40120 & T_4329_43;
  assign T_40122 = T_40121 & T_4329_42;
  assign T_40123 = T_40122 & T_4329_41;
  assign T_40139 = T_39738 & T_4334_45;
  assign T_40140 = T_40139 & T_4334_44;
  assign T_40141 = T_40140 & T_4334_43;
  assign T_40142 = T_40141 & T_4334_42;
  assign T_40143 = T_40142 & T_4334_41;
  assign T_40158 = T_39677 & T_4319_46;
  assign T_40159 = T_40158 & T_4319_45;
  assign T_40160 = T_40159 & T_4319_44;
  assign T_40161 = T_40160 & T_4319_43;
  assign T_40162 = T_40161 & T_4319_42;
  assign T_40163 = T_40162 & T_4319_41;
  assign T_40178 = T_39697 & T_4324_46;
  assign T_40179 = T_40178 & T_4324_45;
  assign T_40180 = T_40179 & T_4324_44;
  assign T_40181 = T_40180 & T_4324_43;
  assign T_40182 = T_40181 & T_4324_42;
  assign T_40183 = T_40182 & T_4324_41;
  assign T_40198 = T_39717 & T_4329_46;
  assign T_40199 = T_40198 & T_4329_45;
  assign T_40200 = T_40199 & T_4329_44;
  assign T_40201 = T_40200 & T_4329_43;
  assign T_40202 = T_40201 & T_4329_42;
  assign T_40203 = T_40202 & T_4329_41;
  assign T_40218 = T_39737 & T_4334_46;
  assign T_40219 = T_40218 & T_4334_45;
  assign T_40220 = T_40219 & T_4334_44;
  assign T_40221 = T_40220 & T_4334_43;
  assign T_40222 = T_40221 & T_4334_42;
  assign T_40223 = T_40222 & T_4334_41;
  assign T_40237 = T_39676 & T_4319_47;
  assign T_40238 = T_40237 & T_4319_46;
  assign T_40239 = T_40238 & T_4319_45;
  assign T_40240 = T_40239 & T_4319_44;
  assign T_40241 = T_40240 & T_4319_43;
  assign T_40242 = T_40241 & T_4319_42;
  assign T_40243 = T_40242 & T_4319_41;
  assign T_40257 = T_39696 & T_4324_47;
  assign T_40258 = T_40257 & T_4324_46;
  assign T_40259 = T_40258 & T_4324_45;
  assign T_40260 = T_40259 & T_4324_44;
  assign T_40261 = T_40260 & T_4324_43;
  assign T_40262 = T_40261 & T_4324_42;
  assign T_40263 = T_40262 & T_4324_41;
  assign T_40277 = T_39716 & T_4329_47;
  assign T_40278 = T_40277 & T_4329_46;
  assign T_40279 = T_40278 & T_4329_45;
  assign T_40280 = T_40279 & T_4329_44;
  assign T_40281 = T_40280 & T_4329_43;
  assign T_40282 = T_40281 & T_4329_42;
  assign T_40283 = T_40282 & T_4329_41;
  assign T_40297 = T_39736 & T_4334_47;
  assign T_40298 = T_40297 & T_4334_46;
  assign T_40299 = T_40298 & T_4334_45;
  assign T_40300 = T_40299 & T_4334_44;
  assign T_40301 = T_40300 & T_4334_43;
  assign T_40302 = T_40301 & T_4334_42;
  assign T_40303 = T_40302 & T_4334_41;
  assign T_40316 = T_39675 & T_4319_48;
  assign T_40317 = T_40316 & T_4319_47;
  assign T_40318 = T_40317 & T_4319_46;
  assign T_40319 = T_40318 & T_4319_45;
  assign T_40320 = T_40319 & T_4319_44;
  assign T_40321 = T_40320 & T_4319_43;
  assign T_40322 = T_40321 & T_4319_42;
  assign T_40323 = T_40322 & T_4319_41;
  assign T_40336 = T_39695 & T_4324_48;
  assign T_40337 = T_40336 & T_4324_47;
  assign T_40338 = T_40337 & T_4324_46;
  assign T_40339 = T_40338 & T_4324_45;
  assign T_40340 = T_40339 & T_4324_44;
  assign T_40341 = T_40340 & T_4324_43;
  assign T_40342 = T_40341 & T_4324_42;
  assign T_40343 = T_40342 & T_4324_41;
  assign T_40356 = T_39715 & T_4329_48;
  assign T_40357 = T_40356 & T_4329_47;
  assign T_40358 = T_40357 & T_4329_46;
  assign T_40359 = T_40358 & T_4329_45;
  assign T_40360 = T_40359 & T_4329_44;
  assign T_40361 = T_40360 & T_4329_43;
  assign T_40362 = T_40361 & T_4329_42;
  assign T_40363 = T_40362 & T_4329_41;
  assign T_40376 = T_39735 & T_4334_48;
  assign T_40377 = T_40376 & T_4334_47;
  assign T_40378 = T_40377 & T_4334_46;
  assign T_40379 = T_40378 & T_4334_45;
  assign T_40380 = T_40379 & T_4334_44;
  assign T_40381 = T_40380 & T_4334_43;
  assign T_40382 = T_40381 & T_4334_42;
  assign T_40383 = T_40382 & T_4334_41;
  assign T_40395 = T_39674 & T_4319_49;
  assign T_40396 = T_40395 & T_4319_48;
  assign T_40397 = T_40396 & T_4319_47;
  assign T_40398 = T_40397 & T_4319_46;
  assign T_40399 = T_40398 & T_4319_45;
  assign T_40400 = T_40399 & T_4319_44;
  assign T_40401 = T_40400 & T_4319_43;
  assign T_40402 = T_40401 & T_4319_42;
  assign T_40403 = T_40402 & T_4319_41;
  assign T_40415 = T_39694 & T_4324_49;
  assign T_40416 = T_40415 & T_4324_48;
  assign T_40417 = T_40416 & T_4324_47;
  assign T_40418 = T_40417 & T_4324_46;
  assign T_40419 = T_40418 & T_4324_45;
  assign T_40420 = T_40419 & T_4324_44;
  assign T_40421 = T_40420 & T_4324_43;
  assign T_40422 = T_40421 & T_4324_42;
  assign T_40423 = T_40422 & T_4324_41;
  assign T_40435 = T_39714 & T_4329_49;
  assign T_40436 = T_40435 & T_4329_48;
  assign T_40437 = T_40436 & T_4329_47;
  assign T_40438 = T_40437 & T_4329_46;
  assign T_40439 = T_40438 & T_4329_45;
  assign T_40440 = T_40439 & T_4329_44;
  assign T_40441 = T_40440 & T_4329_43;
  assign T_40442 = T_40441 & T_4329_42;
  assign T_40443 = T_40442 & T_4329_41;
  assign T_40455 = T_39734 & T_4334_49;
  assign T_40456 = T_40455 & T_4334_48;
  assign T_40457 = T_40456 & T_4334_47;
  assign T_40458 = T_40457 & T_4334_46;
  assign T_40459 = T_40458 & T_4334_45;
  assign T_40460 = T_40459 & T_4334_44;
  assign T_40461 = T_40460 & T_4334_43;
  assign T_40462 = T_40461 & T_4334_42;
  assign T_40463 = T_40462 & T_4334_41;
  assign T_40474 = T_39673 & T_4319_50;
  assign T_40475 = T_40474 & T_4319_49;
  assign T_40476 = T_40475 & T_4319_48;
  assign T_40477 = T_40476 & T_4319_47;
  assign T_40478 = T_40477 & T_4319_46;
  assign T_40479 = T_40478 & T_4319_45;
  assign T_40480 = T_40479 & T_4319_44;
  assign T_40481 = T_40480 & T_4319_43;
  assign T_40482 = T_40481 & T_4319_42;
  assign T_40483 = T_40482 & T_4319_41;
  assign T_40494 = T_39693 & T_4324_50;
  assign T_40495 = T_40494 & T_4324_49;
  assign T_40496 = T_40495 & T_4324_48;
  assign T_40497 = T_40496 & T_4324_47;
  assign T_40498 = T_40497 & T_4324_46;
  assign T_40499 = T_40498 & T_4324_45;
  assign T_40500 = T_40499 & T_4324_44;
  assign T_40501 = T_40500 & T_4324_43;
  assign T_40502 = T_40501 & T_4324_42;
  assign T_40503 = T_40502 & T_4324_41;
  assign T_40514 = T_39713 & T_4329_50;
  assign T_40515 = T_40514 & T_4329_49;
  assign T_40516 = T_40515 & T_4329_48;
  assign T_40517 = T_40516 & T_4329_47;
  assign T_40518 = T_40517 & T_4329_46;
  assign T_40519 = T_40518 & T_4329_45;
  assign T_40520 = T_40519 & T_4329_44;
  assign T_40521 = T_40520 & T_4329_43;
  assign T_40522 = T_40521 & T_4329_42;
  assign T_40523 = T_40522 & T_4329_41;
  assign T_40534 = T_39733 & T_4334_50;
  assign T_40535 = T_40534 & T_4334_49;
  assign T_40536 = T_40535 & T_4334_48;
  assign T_40537 = T_40536 & T_4334_47;
  assign T_40538 = T_40537 & T_4334_46;
  assign T_40539 = T_40538 & T_4334_45;
  assign T_40540 = T_40539 & T_4334_44;
  assign T_40541 = T_40540 & T_4334_43;
  assign T_40542 = T_40541 & T_4334_42;
  assign T_40543 = T_40542 & T_4334_41;
  assign T_40553 = T_39672 & T_4319_51;
  assign T_40554 = T_40553 & T_4319_50;
  assign T_40555 = T_40554 & T_4319_49;
  assign T_40556 = T_40555 & T_4319_48;
  assign T_40557 = T_40556 & T_4319_47;
  assign T_40558 = T_40557 & T_4319_46;
  assign T_40559 = T_40558 & T_4319_45;
  assign T_40560 = T_40559 & T_4319_44;
  assign T_40561 = T_40560 & T_4319_43;
  assign T_40562 = T_40561 & T_4319_42;
  assign T_40563 = T_40562 & T_4319_41;
  assign T_40573 = T_39692 & T_4324_51;
  assign T_40574 = T_40573 & T_4324_50;
  assign T_40575 = T_40574 & T_4324_49;
  assign T_40576 = T_40575 & T_4324_48;
  assign T_40577 = T_40576 & T_4324_47;
  assign T_40578 = T_40577 & T_4324_46;
  assign T_40579 = T_40578 & T_4324_45;
  assign T_40580 = T_40579 & T_4324_44;
  assign T_40581 = T_40580 & T_4324_43;
  assign T_40582 = T_40581 & T_4324_42;
  assign T_40583 = T_40582 & T_4324_41;
  assign T_40593 = T_39712 & T_4329_51;
  assign T_40594 = T_40593 & T_4329_50;
  assign T_40595 = T_40594 & T_4329_49;
  assign T_40596 = T_40595 & T_4329_48;
  assign T_40597 = T_40596 & T_4329_47;
  assign T_40598 = T_40597 & T_4329_46;
  assign T_40599 = T_40598 & T_4329_45;
  assign T_40600 = T_40599 & T_4329_44;
  assign T_40601 = T_40600 & T_4329_43;
  assign T_40602 = T_40601 & T_4329_42;
  assign T_40603 = T_40602 & T_4329_41;
  assign T_40613 = T_39732 & T_4334_51;
  assign T_40614 = T_40613 & T_4334_50;
  assign T_40615 = T_40614 & T_4334_49;
  assign T_40616 = T_40615 & T_4334_48;
  assign T_40617 = T_40616 & T_4334_47;
  assign T_40618 = T_40617 & T_4334_46;
  assign T_40619 = T_40618 & T_4334_45;
  assign T_40620 = T_40619 & T_4334_44;
  assign T_40621 = T_40620 & T_4334_43;
  assign T_40622 = T_40621 & T_4334_42;
  assign T_40623 = T_40622 & T_4334_41;
  assign T_40632 = T_39671 & T_4319_52;
  assign T_40633 = T_40632 & T_4319_51;
  assign T_40634 = T_40633 & T_4319_50;
  assign T_40635 = T_40634 & T_4319_49;
  assign T_40636 = T_40635 & T_4319_48;
  assign T_40637 = T_40636 & T_4319_47;
  assign T_40638 = T_40637 & T_4319_46;
  assign T_40639 = T_40638 & T_4319_45;
  assign T_40640 = T_40639 & T_4319_44;
  assign T_40641 = T_40640 & T_4319_43;
  assign T_40642 = T_40641 & T_4319_42;
  assign T_40643 = T_40642 & T_4319_41;
  assign T_40652 = T_39691 & T_4324_52;
  assign T_40653 = T_40652 & T_4324_51;
  assign T_40654 = T_40653 & T_4324_50;
  assign T_40655 = T_40654 & T_4324_49;
  assign T_40656 = T_40655 & T_4324_48;
  assign T_40657 = T_40656 & T_4324_47;
  assign T_40658 = T_40657 & T_4324_46;
  assign T_40659 = T_40658 & T_4324_45;
  assign T_40660 = T_40659 & T_4324_44;
  assign T_40661 = T_40660 & T_4324_43;
  assign T_40662 = T_40661 & T_4324_42;
  assign T_40663 = T_40662 & T_4324_41;
  assign T_40672 = T_39711 & T_4329_52;
  assign T_40673 = T_40672 & T_4329_51;
  assign T_40674 = T_40673 & T_4329_50;
  assign T_40675 = T_40674 & T_4329_49;
  assign T_40676 = T_40675 & T_4329_48;
  assign T_40677 = T_40676 & T_4329_47;
  assign T_40678 = T_40677 & T_4329_46;
  assign T_40679 = T_40678 & T_4329_45;
  assign T_40680 = T_40679 & T_4329_44;
  assign T_40681 = T_40680 & T_4329_43;
  assign T_40682 = T_40681 & T_4329_42;
  assign T_40683 = T_40682 & T_4329_41;
  assign T_40692 = T_39731 & T_4334_52;
  assign T_40693 = T_40692 & T_4334_51;
  assign T_40694 = T_40693 & T_4334_50;
  assign T_40695 = T_40694 & T_4334_49;
  assign T_40696 = T_40695 & T_4334_48;
  assign T_40697 = T_40696 & T_4334_47;
  assign T_40698 = T_40697 & T_4334_46;
  assign T_40699 = T_40698 & T_4334_45;
  assign T_40700 = T_40699 & T_4334_44;
  assign T_40701 = T_40700 & T_4334_43;
  assign T_40702 = T_40701 & T_4334_42;
  assign T_40703 = T_40702 & T_4334_41;
  assign T_40711 = T_39670 & T_4319_53;
  assign T_40712 = T_40711 & T_4319_52;
  assign T_40713 = T_40712 & T_4319_51;
  assign T_40714 = T_40713 & T_4319_50;
  assign T_40715 = T_40714 & T_4319_49;
  assign T_40716 = T_40715 & T_4319_48;
  assign T_40717 = T_40716 & T_4319_47;
  assign T_40718 = T_40717 & T_4319_46;
  assign T_40719 = T_40718 & T_4319_45;
  assign T_40720 = T_40719 & T_4319_44;
  assign T_40721 = T_40720 & T_4319_43;
  assign T_40722 = T_40721 & T_4319_42;
  assign T_40723 = T_40722 & T_4319_41;
  assign T_40731 = T_39690 & T_4324_53;
  assign T_40732 = T_40731 & T_4324_52;
  assign T_40733 = T_40732 & T_4324_51;
  assign T_40734 = T_40733 & T_4324_50;
  assign T_40735 = T_40734 & T_4324_49;
  assign T_40736 = T_40735 & T_4324_48;
  assign T_40737 = T_40736 & T_4324_47;
  assign T_40738 = T_40737 & T_4324_46;
  assign T_40739 = T_40738 & T_4324_45;
  assign T_40740 = T_40739 & T_4324_44;
  assign T_40741 = T_40740 & T_4324_43;
  assign T_40742 = T_40741 & T_4324_42;
  assign T_40743 = T_40742 & T_4324_41;
  assign T_40751 = T_39710 & T_4329_53;
  assign T_40752 = T_40751 & T_4329_52;
  assign T_40753 = T_40752 & T_4329_51;
  assign T_40754 = T_40753 & T_4329_50;
  assign T_40755 = T_40754 & T_4329_49;
  assign T_40756 = T_40755 & T_4329_48;
  assign T_40757 = T_40756 & T_4329_47;
  assign T_40758 = T_40757 & T_4329_46;
  assign T_40759 = T_40758 & T_4329_45;
  assign T_40760 = T_40759 & T_4329_44;
  assign T_40761 = T_40760 & T_4329_43;
  assign T_40762 = T_40761 & T_4329_42;
  assign T_40763 = T_40762 & T_4329_41;
  assign T_40771 = T_39730 & T_4334_53;
  assign T_40772 = T_40771 & T_4334_52;
  assign T_40773 = T_40772 & T_4334_51;
  assign T_40774 = T_40773 & T_4334_50;
  assign T_40775 = T_40774 & T_4334_49;
  assign T_40776 = T_40775 & T_4334_48;
  assign T_40777 = T_40776 & T_4334_47;
  assign T_40778 = T_40777 & T_4334_46;
  assign T_40779 = T_40778 & T_4334_45;
  assign T_40780 = T_40779 & T_4334_44;
  assign T_40781 = T_40780 & T_4334_43;
  assign T_40782 = T_40781 & T_4334_42;
  assign T_40783 = T_40782 & T_4334_41;
  assign T_40790 = T_39669 & T_4319_54;
  assign T_40791 = T_40790 & T_4319_53;
  assign T_40792 = T_40791 & T_4319_52;
  assign T_40793 = T_40792 & T_4319_51;
  assign T_40794 = T_40793 & T_4319_50;
  assign T_40795 = T_40794 & T_4319_49;
  assign T_40796 = T_40795 & T_4319_48;
  assign T_40797 = T_40796 & T_4319_47;
  assign T_40798 = T_40797 & T_4319_46;
  assign T_40799 = T_40798 & T_4319_45;
  assign T_40800 = T_40799 & T_4319_44;
  assign T_40801 = T_40800 & T_4319_43;
  assign T_40802 = T_40801 & T_4319_42;
  assign T_40803 = T_40802 & T_4319_41;
  assign T_40810 = T_39689 & T_4324_54;
  assign T_40811 = T_40810 & T_4324_53;
  assign T_40812 = T_40811 & T_4324_52;
  assign T_40813 = T_40812 & T_4324_51;
  assign T_40814 = T_40813 & T_4324_50;
  assign T_40815 = T_40814 & T_4324_49;
  assign T_40816 = T_40815 & T_4324_48;
  assign T_40817 = T_40816 & T_4324_47;
  assign T_40818 = T_40817 & T_4324_46;
  assign T_40819 = T_40818 & T_4324_45;
  assign T_40820 = T_40819 & T_4324_44;
  assign T_40821 = T_40820 & T_4324_43;
  assign T_40822 = T_40821 & T_4324_42;
  assign T_40823 = T_40822 & T_4324_41;
  assign T_40830 = T_39709 & T_4329_54;
  assign T_40831 = T_40830 & T_4329_53;
  assign T_40832 = T_40831 & T_4329_52;
  assign T_40833 = T_40832 & T_4329_51;
  assign T_40834 = T_40833 & T_4329_50;
  assign T_40835 = T_40834 & T_4329_49;
  assign T_40836 = T_40835 & T_4329_48;
  assign T_40837 = T_40836 & T_4329_47;
  assign T_40838 = T_40837 & T_4329_46;
  assign T_40839 = T_40838 & T_4329_45;
  assign T_40840 = T_40839 & T_4329_44;
  assign T_40841 = T_40840 & T_4329_43;
  assign T_40842 = T_40841 & T_4329_42;
  assign T_40843 = T_40842 & T_4329_41;
  assign T_40850 = T_39729 & T_4334_54;
  assign T_40851 = T_40850 & T_4334_53;
  assign T_40852 = T_40851 & T_4334_52;
  assign T_40853 = T_40852 & T_4334_51;
  assign T_40854 = T_40853 & T_4334_50;
  assign T_40855 = T_40854 & T_4334_49;
  assign T_40856 = T_40855 & T_4334_48;
  assign T_40857 = T_40856 & T_4334_47;
  assign T_40858 = T_40857 & T_4334_46;
  assign T_40859 = T_40858 & T_4334_45;
  assign T_40860 = T_40859 & T_4334_44;
  assign T_40861 = T_40860 & T_4334_43;
  assign T_40862 = T_40861 & T_4334_42;
  assign T_40863 = T_40862 & T_4334_41;
  assign T_40869 = T_39668 & T_4319_55;
  assign T_40870 = T_40869 & T_4319_54;
  assign T_40871 = T_40870 & T_4319_53;
  assign T_40872 = T_40871 & T_4319_52;
  assign T_40873 = T_40872 & T_4319_51;
  assign T_40874 = T_40873 & T_4319_50;
  assign T_40875 = T_40874 & T_4319_49;
  assign T_40876 = T_40875 & T_4319_48;
  assign T_40877 = T_40876 & T_4319_47;
  assign T_40878 = T_40877 & T_4319_46;
  assign T_40879 = T_40878 & T_4319_45;
  assign T_40880 = T_40879 & T_4319_44;
  assign T_40881 = T_40880 & T_4319_43;
  assign T_40882 = T_40881 & T_4319_42;
  assign T_40883 = T_40882 & T_4319_41;
  assign T_40889 = T_39688 & T_4324_55;
  assign T_40890 = T_40889 & T_4324_54;
  assign T_40891 = T_40890 & T_4324_53;
  assign T_40892 = T_40891 & T_4324_52;
  assign T_40893 = T_40892 & T_4324_51;
  assign T_40894 = T_40893 & T_4324_50;
  assign T_40895 = T_40894 & T_4324_49;
  assign T_40896 = T_40895 & T_4324_48;
  assign T_40897 = T_40896 & T_4324_47;
  assign T_40898 = T_40897 & T_4324_46;
  assign T_40899 = T_40898 & T_4324_45;
  assign T_40900 = T_40899 & T_4324_44;
  assign T_40901 = T_40900 & T_4324_43;
  assign T_40902 = T_40901 & T_4324_42;
  assign T_40903 = T_40902 & T_4324_41;
  assign T_40909 = T_39708 & T_4329_55;
  assign T_40910 = T_40909 & T_4329_54;
  assign T_40911 = T_40910 & T_4329_53;
  assign T_40912 = T_40911 & T_4329_52;
  assign T_40913 = T_40912 & T_4329_51;
  assign T_40914 = T_40913 & T_4329_50;
  assign T_40915 = T_40914 & T_4329_49;
  assign T_40916 = T_40915 & T_4329_48;
  assign T_40917 = T_40916 & T_4329_47;
  assign T_40918 = T_40917 & T_4329_46;
  assign T_40919 = T_40918 & T_4329_45;
  assign T_40920 = T_40919 & T_4329_44;
  assign T_40921 = T_40920 & T_4329_43;
  assign T_40922 = T_40921 & T_4329_42;
  assign T_40923 = T_40922 & T_4329_41;
  assign T_40929 = T_39728 & T_4334_55;
  assign T_40930 = T_40929 & T_4334_54;
  assign T_40931 = T_40930 & T_4334_53;
  assign T_40932 = T_40931 & T_4334_52;
  assign T_40933 = T_40932 & T_4334_51;
  assign T_40934 = T_40933 & T_4334_50;
  assign T_40935 = T_40934 & T_4334_49;
  assign T_40936 = T_40935 & T_4334_48;
  assign T_40937 = T_40936 & T_4334_47;
  assign T_40938 = T_40937 & T_4334_46;
  assign T_40939 = T_40938 & T_4334_45;
  assign T_40940 = T_40939 & T_4334_44;
  assign T_40941 = T_40940 & T_4334_43;
  assign T_40942 = T_40941 & T_4334_42;
  assign T_40943 = T_40942 & T_4334_41;
  assign T_40948 = T_39667 & T_4319_56;
  assign T_40949 = T_40948 & T_4319_55;
  assign T_40950 = T_40949 & T_4319_54;
  assign T_40951 = T_40950 & T_4319_53;
  assign T_40952 = T_40951 & T_4319_52;
  assign T_40953 = T_40952 & T_4319_51;
  assign T_40954 = T_40953 & T_4319_50;
  assign T_40955 = T_40954 & T_4319_49;
  assign T_40956 = T_40955 & T_4319_48;
  assign T_40957 = T_40956 & T_4319_47;
  assign T_40958 = T_40957 & T_4319_46;
  assign T_40959 = T_40958 & T_4319_45;
  assign T_40960 = T_40959 & T_4319_44;
  assign T_40961 = T_40960 & T_4319_43;
  assign T_40962 = T_40961 & T_4319_42;
  assign T_40963 = T_40962 & T_4319_41;
  assign T_40968 = T_39687 & T_4324_56;
  assign T_40969 = T_40968 & T_4324_55;
  assign T_40970 = T_40969 & T_4324_54;
  assign T_40971 = T_40970 & T_4324_53;
  assign T_40972 = T_40971 & T_4324_52;
  assign T_40973 = T_40972 & T_4324_51;
  assign T_40974 = T_40973 & T_4324_50;
  assign T_40975 = T_40974 & T_4324_49;
  assign T_40976 = T_40975 & T_4324_48;
  assign T_40977 = T_40976 & T_4324_47;
  assign T_40978 = T_40977 & T_4324_46;
  assign T_40979 = T_40978 & T_4324_45;
  assign T_40980 = T_40979 & T_4324_44;
  assign T_40981 = T_40980 & T_4324_43;
  assign T_40982 = T_40981 & T_4324_42;
  assign T_40983 = T_40982 & T_4324_41;
  assign T_40988 = T_39707 & T_4329_56;
  assign T_40989 = T_40988 & T_4329_55;
  assign T_40990 = T_40989 & T_4329_54;
  assign T_40991 = T_40990 & T_4329_53;
  assign T_40992 = T_40991 & T_4329_52;
  assign T_40993 = T_40992 & T_4329_51;
  assign T_40994 = T_40993 & T_4329_50;
  assign T_40995 = T_40994 & T_4329_49;
  assign T_40996 = T_40995 & T_4329_48;
  assign T_40997 = T_40996 & T_4329_47;
  assign T_40998 = T_40997 & T_4329_46;
  assign T_40999 = T_40998 & T_4329_45;
  assign T_41000 = T_40999 & T_4329_44;
  assign T_41001 = T_41000 & T_4329_43;
  assign T_41002 = T_41001 & T_4329_42;
  assign T_41003 = T_41002 & T_4329_41;
  assign T_41008 = T_39727 & T_4334_56;
  assign T_41009 = T_41008 & T_4334_55;
  assign T_41010 = T_41009 & T_4334_54;
  assign T_41011 = T_41010 & T_4334_53;
  assign T_41012 = T_41011 & T_4334_52;
  assign T_41013 = T_41012 & T_4334_51;
  assign T_41014 = T_41013 & T_4334_50;
  assign T_41015 = T_41014 & T_4334_49;
  assign T_41016 = T_41015 & T_4334_48;
  assign T_41017 = T_41016 & T_4334_47;
  assign T_41018 = T_41017 & T_4334_46;
  assign T_41019 = T_41018 & T_4334_45;
  assign T_41020 = T_41019 & T_4334_44;
  assign T_41021 = T_41020 & T_4334_43;
  assign T_41022 = T_41021 & T_4334_42;
  assign T_41023 = T_41022 & T_4334_41;
  assign T_41027 = T_39666 & T_4319_57;
  assign T_41028 = T_41027 & T_4319_56;
  assign T_41029 = T_41028 & T_4319_55;
  assign T_41030 = T_41029 & T_4319_54;
  assign T_41031 = T_41030 & T_4319_53;
  assign T_41032 = T_41031 & T_4319_52;
  assign T_41033 = T_41032 & T_4319_51;
  assign T_41034 = T_41033 & T_4319_50;
  assign T_41035 = T_41034 & T_4319_49;
  assign T_41036 = T_41035 & T_4319_48;
  assign T_41037 = T_41036 & T_4319_47;
  assign T_41038 = T_41037 & T_4319_46;
  assign T_41039 = T_41038 & T_4319_45;
  assign T_41040 = T_41039 & T_4319_44;
  assign T_41041 = T_41040 & T_4319_43;
  assign T_41042 = T_41041 & T_4319_42;
  assign T_41043 = T_41042 & T_4319_41;
  assign T_41047 = T_39686 & T_4324_57;
  assign T_41048 = T_41047 & T_4324_56;
  assign T_41049 = T_41048 & T_4324_55;
  assign T_41050 = T_41049 & T_4324_54;
  assign T_41051 = T_41050 & T_4324_53;
  assign T_41052 = T_41051 & T_4324_52;
  assign T_41053 = T_41052 & T_4324_51;
  assign T_41054 = T_41053 & T_4324_50;
  assign T_41055 = T_41054 & T_4324_49;
  assign T_41056 = T_41055 & T_4324_48;
  assign T_41057 = T_41056 & T_4324_47;
  assign T_41058 = T_41057 & T_4324_46;
  assign T_41059 = T_41058 & T_4324_45;
  assign T_41060 = T_41059 & T_4324_44;
  assign T_41061 = T_41060 & T_4324_43;
  assign T_41062 = T_41061 & T_4324_42;
  assign T_41063 = T_41062 & T_4324_41;
  assign T_41067 = T_39706 & T_4329_57;
  assign T_41068 = T_41067 & T_4329_56;
  assign T_41069 = T_41068 & T_4329_55;
  assign T_41070 = T_41069 & T_4329_54;
  assign T_41071 = T_41070 & T_4329_53;
  assign T_41072 = T_41071 & T_4329_52;
  assign T_41073 = T_41072 & T_4329_51;
  assign T_41074 = T_41073 & T_4329_50;
  assign T_41075 = T_41074 & T_4329_49;
  assign T_41076 = T_41075 & T_4329_48;
  assign T_41077 = T_41076 & T_4329_47;
  assign T_41078 = T_41077 & T_4329_46;
  assign T_41079 = T_41078 & T_4329_45;
  assign T_41080 = T_41079 & T_4329_44;
  assign T_41081 = T_41080 & T_4329_43;
  assign T_41082 = T_41081 & T_4329_42;
  assign T_41083 = T_41082 & T_4329_41;
  assign T_41087 = T_39726 & T_4334_57;
  assign T_41088 = T_41087 & T_4334_56;
  assign T_41089 = T_41088 & T_4334_55;
  assign T_41090 = T_41089 & T_4334_54;
  assign T_41091 = T_41090 & T_4334_53;
  assign T_41092 = T_41091 & T_4334_52;
  assign T_41093 = T_41092 & T_4334_51;
  assign T_41094 = T_41093 & T_4334_50;
  assign T_41095 = T_41094 & T_4334_49;
  assign T_41096 = T_41095 & T_4334_48;
  assign T_41097 = T_41096 & T_4334_47;
  assign T_41098 = T_41097 & T_4334_46;
  assign T_41099 = T_41098 & T_4334_45;
  assign T_41100 = T_41099 & T_4334_44;
  assign T_41101 = T_41100 & T_4334_43;
  assign T_41102 = T_41101 & T_4334_42;
  assign T_41103 = T_41102 & T_4334_41;
  assign T_41106 = T_39665 & T_4319_58;
  assign T_41107 = T_41106 & T_4319_57;
  assign T_41108 = T_41107 & T_4319_56;
  assign T_41109 = T_41108 & T_4319_55;
  assign T_41110 = T_41109 & T_4319_54;
  assign T_41111 = T_41110 & T_4319_53;
  assign T_41112 = T_41111 & T_4319_52;
  assign T_41113 = T_41112 & T_4319_51;
  assign T_41114 = T_41113 & T_4319_50;
  assign T_41115 = T_41114 & T_4319_49;
  assign T_41116 = T_41115 & T_4319_48;
  assign T_41117 = T_41116 & T_4319_47;
  assign T_41118 = T_41117 & T_4319_46;
  assign T_41119 = T_41118 & T_4319_45;
  assign T_41120 = T_41119 & T_4319_44;
  assign T_41121 = T_41120 & T_4319_43;
  assign T_41122 = T_41121 & T_4319_42;
  assign T_41123 = T_41122 & T_4319_41;
  assign T_41126 = T_39685 & T_4324_58;
  assign T_41127 = T_41126 & T_4324_57;
  assign T_41128 = T_41127 & T_4324_56;
  assign T_41129 = T_41128 & T_4324_55;
  assign T_41130 = T_41129 & T_4324_54;
  assign T_41131 = T_41130 & T_4324_53;
  assign T_41132 = T_41131 & T_4324_52;
  assign T_41133 = T_41132 & T_4324_51;
  assign T_41134 = T_41133 & T_4324_50;
  assign T_41135 = T_41134 & T_4324_49;
  assign T_41136 = T_41135 & T_4324_48;
  assign T_41137 = T_41136 & T_4324_47;
  assign T_41138 = T_41137 & T_4324_46;
  assign T_41139 = T_41138 & T_4324_45;
  assign T_41140 = T_41139 & T_4324_44;
  assign T_41141 = T_41140 & T_4324_43;
  assign T_41142 = T_41141 & T_4324_42;
  assign T_41143 = T_41142 & T_4324_41;
  assign T_41146 = T_39705 & T_4329_58;
  assign T_41147 = T_41146 & T_4329_57;
  assign T_41148 = T_41147 & T_4329_56;
  assign T_41149 = T_41148 & T_4329_55;
  assign T_41150 = T_41149 & T_4329_54;
  assign T_41151 = T_41150 & T_4329_53;
  assign T_41152 = T_41151 & T_4329_52;
  assign T_41153 = T_41152 & T_4329_51;
  assign T_41154 = T_41153 & T_4329_50;
  assign T_41155 = T_41154 & T_4329_49;
  assign T_41156 = T_41155 & T_4329_48;
  assign T_41157 = T_41156 & T_4329_47;
  assign T_41158 = T_41157 & T_4329_46;
  assign T_41159 = T_41158 & T_4329_45;
  assign T_41160 = T_41159 & T_4329_44;
  assign T_41161 = T_41160 & T_4329_43;
  assign T_41162 = T_41161 & T_4329_42;
  assign T_41163 = T_41162 & T_4329_41;
  assign T_41166 = T_39725 & T_4334_58;
  assign T_41167 = T_41166 & T_4334_57;
  assign T_41168 = T_41167 & T_4334_56;
  assign T_41169 = T_41168 & T_4334_55;
  assign T_41170 = T_41169 & T_4334_54;
  assign T_41171 = T_41170 & T_4334_53;
  assign T_41172 = T_41171 & T_4334_52;
  assign T_41173 = T_41172 & T_4334_51;
  assign T_41174 = T_41173 & T_4334_50;
  assign T_41175 = T_41174 & T_4334_49;
  assign T_41176 = T_41175 & T_4334_48;
  assign T_41177 = T_41176 & T_4334_47;
  assign T_41178 = T_41177 & T_4334_46;
  assign T_41179 = T_41178 & T_4334_45;
  assign T_41180 = T_41179 & T_4334_44;
  assign T_41181 = T_41180 & T_4334_43;
  assign T_41182 = T_41181 & T_4334_42;
  assign T_41183 = T_41182 & T_4334_41;
  assign T_41185 = T_27876 & T_4319_59;
  assign T_41186 = T_41185 & T_4319_58;
  assign T_41187 = T_41186 & T_4319_57;
  assign T_41188 = T_41187 & T_4319_56;
  assign T_41189 = T_41188 & T_4319_55;
  assign T_41190 = T_41189 & T_4319_54;
  assign T_41191 = T_41190 & T_4319_53;
  assign T_41192 = T_41191 & T_4319_52;
  assign T_41193 = T_41192 & T_4319_51;
  assign T_41194 = T_41193 & T_4319_50;
  assign T_41195 = T_41194 & T_4319_49;
  assign T_41196 = T_41195 & T_4319_48;
  assign T_41197 = T_41196 & T_4319_47;
  assign T_41198 = T_41197 & T_4319_46;
  assign T_41199 = T_41198 & T_4319_45;
  assign T_41200 = T_41199 & T_4319_44;
  assign T_41201 = T_41200 & T_4319_43;
  assign T_41202 = T_41201 & T_4319_42;
  assign T_41203 = T_41202 & T_4319_41;
  assign T_41205 = T_27882 & T_4324_59;
  assign T_41206 = T_41205 & T_4324_58;
  assign T_41207 = T_41206 & T_4324_57;
  assign T_41208 = T_41207 & T_4324_56;
  assign T_41209 = T_41208 & T_4324_55;
  assign T_41210 = T_41209 & T_4324_54;
  assign T_41211 = T_41210 & T_4324_53;
  assign T_41212 = T_41211 & T_4324_52;
  assign T_41213 = T_41212 & T_4324_51;
  assign T_41214 = T_41213 & T_4324_50;
  assign T_41215 = T_41214 & T_4324_49;
  assign T_41216 = T_41215 & T_4324_48;
  assign T_41217 = T_41216 & T_4324_47;
  assign T_41218 = T_41217 & T_4324_46;
  assign T_41219 = T_41218 & T_4324_45;
  assign T_41220 = T_41219 & T_4324_44;
  assign T_41221 = T_41220 & T_4324_43;
  assign T_41222 = T_41221 & T_4324_42;
  assign T_41223 = T_41222 & T_4324_41;
  assign T_41225 = T_27886 & T_4329_59;
  assign T_41226 = T_41225 & T_4329_58;
  assign T_41227 = T_41226 & T_4329_57;
  assign T_41228 = T_41227 & T_4329_56;
  assign T_41229 = T_41228 & T_4329_55;
  assign T_41230 = T_41229 & T_4329_54;
  assign T_41231 = T_41230 & T_4329_53;
  assign T_41232 = T_41231 & T_4329_52;
  assign T_41233 = T_41232 & T_4329_51;
  assign T_41234 = T_41233 & T_4329_50;
  assign T_41235 = T_41234 & T_4329_49;
  assign T_41236 = T_41235 & T_4329_48;
  assign T_41237 = T_41236 & T_4329_47;
  assign T_41238 = T_41237 & T_4329_46;
  assign T_41239 = T_41238 & T_4329_45;
  assign T_41240 = T_41239 & T_4329_44;
  assign T_41241 = T_41240 & T_4329_43;
  assign T_41242 = T_41241 & T_4329_42;
  assign T_41243 = T_41242 & T_4329_41;
  assign T_41245 = T_27892 & T_4334_59;
  assign T_41246 = T_41245 & T_4334_58;
  assign T_41247 = T_41246 & T_4334_57;
  assign T_41248 = T_41247 & T_4334_56;
  assign T_41249 = T_41248 & T_4334_55;
  assign T_41250 = T_41249 & T_4334_54;
  assign T_41251 = T_41250 & T_4334_53;
  assign T_41252 = T_41251 & T_4334_52;
  assign T_41253 = T_41252 & T_4334_51;
  assign T_41254 = T_41253 & T_4334_50;
  assign T_41255 = T_41254 & T_4334_49;
  assign T_41256 = T_41255 & T_4334_48;
  assign T_41257 = T_41256 & T_4334_47;
  assign T_41258 = T_41257 & T_4334_46;
  assign T_41259 = T_41258 & T_4334_45;
  assign T_41260 = T_41259 & T_4334_44;
  assign T_41261 = T_41260 & T_4334_43;
  assign T_41262 = T_41261 & T_4334_42;
  assign T_41263 = T_41262 & T_4334_41;
  assign T_41337 = T_27856 & T_4319_110;
  assign T_41338 = T_41337 & T_4319_109;
  assign T_41339 = T_41338 & T_4319_108;
  assign T_41340 = T_41339 & T_4319_107;
  assign T_41341 = T_41340 & T_4319_106;
  assign T_41342 = T_41341 & T_4319_105;
  assign T_41343 = T_41342 & T_4319_104;
  assign T_41344 = T_41343 & T_4319_103;
  assign T_41345 = T_41344 & T_4319_102;
  assign T_41346 = T_41345 & T_4319_101;
  assign T_41347 = T_41346 & T_4319_100;
  assign T_41348 = T_41347 & T_4319_99;
  assign T_41349 = T_41348 & T_4319_98;
  assign T_41350 = T_41349 & T_4319_97;
  assign T_41351 = T_41350 & T_4319_96;
  assign T_41352 = T_41351 & T_4319_95;
  assign T_41353 = T_41352 & T_4319_94;
  assign T_41354 = T_41353 & T_4319_93;
  assign T_41355 = T_41354 & T_4319_92;
  assign T_41356 = T_41355 & T_4319_91;
  assign T_41357 = T_41356 & T_4319_90;
  assign T_41358 = T_41357 & T_4319_89;
  assign T_41359 = T_41358 & T_4319_88;
  assign T_41360 = T_41359 & T_4319_87;
  assign T_41361 = T_41360 & T_4319_86;
  assign T_41362 = T_41361 & T_4319_85;
  assign T_41363 = T_41362 & T_4319_84;
  assign T_41364 = T_41363 & T_4319_83;
  assign T_41365 = T_41364 & T_4319_82;
  assign T_41366 = T_41365 & T_4319_81;
  assign T_41367 = T_41366 & T_4319_80;
  assign T_41369 = T_27862 & T_4324_110;
  assign T_41370 = T_41369 & T_4324_109;
  assign T_41371 = T_41370 & T_4324_108;
  assign T_41372 = T_41371 & T_4324_107;
  assign T_41373 = T_41372 & T_4324_106;
  assign T_41374 = T_41373 & T_4324_105;
  assign T_41375 = T_41374 & T_4324_104;
  assign T_41376 = T_41375 & T_4324_103;
  assign T_41377 = T_41376 & T_4324_102;
  assign T_41378 = T_41377 & T_4324_101;
  assign T_41379 = T_41378 & T_4324_100;
  assign T_41380 = T_41379 & T_4324_99;
  assign T_41381 = T_41380 & T_4324_98;
  assign T_41382 = T_41381 & T_4324_97;
  assign T_41383 = T_41382 & T_4324_96;
  assign T_41384 = T_41383 & T_4324_95;
  assign T_41385 = T_41384 & T_4324_94;
  assign T_41386 = T_41385 & T_4324_93;
  assign T_41387 = T_41386 & T_4324_92;
  assign T_41388 = T_41387 & T_4324_91;
  assign T_41389 = T_41388 & T_4324_90;
  assign T_41390 = T_41389 & T_4324_89;
  assign T_41391 = T_41390 & T_4324_88;
  assign T_41392 = T_41391 & T_4324_87;
  assign T_41393 = T_41392 & T_4324_86;
  assign T_41394 = T_41393 & T_4324_85;
  assign T_41395 = T_41394 & T_4324_84;
  assign T_41396 = T_41395 & T_4324_83;
  assign T_41397 = T_41396 & T_4324_82;
  assign T_41398 = T_41397 & T_4324_81;
  assign T_41399 = T_41398 & T_4324_80;
  assign T_41401 = T_27866 & T_4329_110;
  assign T_41402 = T_41401 & T_4329_109;
  assign T_41403 = T_41402 & T_4329_108;
  assign T_41404 = T_41403 & T_4329_107;
  assign T_41405 = T_41404 & T_4329_106;
  assign T_41406 = T_41405 & T_4329_105;
  assign T_41407 = T_41406 & T_4329_104;
  assign T_41408 = T_41407 & T_4329_103;
  assign T_41409 = T_41408 & T_4329_102;
  assign T_41410 = T_41409 & T_4329_101;
  assign T_41411 = T_41410 & T_4329_100;
  assign T_41412 = T_41411 & T_4329_99;
  assign T_41413 = T_41412 & T_4329_98;
  assign T_41414 = T_41413 & T_4329_97;
  assign T_41415 = T_41414 & T_4329_96;
  assign T_41416 = T_41415 & T_4329_95;
  assign T_41417 = T_41416 & T_4329_94;
  assign T_41418 = T_41417 & T_4329_93;
  assign T_41419 = T_41418 & T_4329_92;
  assign T_41420 = T_41419 & T_4329_91;
  assign T_41421 = T_41420 & T_4329_90;
  assign T_41422 = T_41421 & T_4329_89;
  assign T_41423 = T_41422 & T_4329_88;
  assign T_41424 = T_41423 & T_4329_87;
  assign T_41425 = T_41424 & T_4329_86;
  assign T_41426 = T_41425 & T_4329_85;
  assign T_41427 = T_41426 & T_4329_84;
  assign T_41428 = T_41427 & T_4329_83;
  assign T_41429 = T_41428 & T_4329_82;
  assign T_41430 = T_41429 & T_4329_81;
  assign T_41431 = T_41430 & T_4329_80;
  assign T_41433 = T_27872 & T_4334_110;
  assign T_41434 = T_41433 & T_4334_109;
  assign T_41435 = T_41434 & T_4334_108;
  assign T_41436 = T_41435 & T_4334_107;
  assign T_41437 = T_41436 & T_4334_106;
  assign T_41438 = T_41437 & T_4334_105;
  assign T_41439 = T_41438 & T_4334_104;
  assign T_41440 = T_41439 & T_4334_103;
  assign T_41441 = T_41440 & T_4334_102;
  assign T_41442 = T_41441 & T_4334_101;
  assign T_41443 = T_41442 & T_4334_100;
  assign T_41444 = T_41443 & T_4334_99;
  assign T_41445 = T_41444 & T_4334_98;
  assign T_41446 = T_41445 & T_4334_97;
  assign T_41447 = T_41446 & T_4334_96;
  assign T_41448 = T_41447 & T_4334_95;
  assign T_41449 = T_41448 & T_4334_94;
  assign T_41450 = T_41449 & T_4334_93;
  assign T_41451 = T_41450 & T_4334_92;
  assign T_41452 = T_41451 & T_4334_91;
  assign T_41453 = T_41452 & T_4334_90;
  assign T_41454 = T_41453 & T_4334_89;
  assign T_41455 = T_41454 & T_4334_88;
  assign T_41456 = T_41455 & T_4334_87;
  assign T_41457 = T_41456 & T_4334_86;
  assign T_41458 = T_41457 & T_4334_85;
  assign T_41459 = T_41458 & T_4334_84;
  assign T_41460 = T_41459 & T_4334_83;
  assign T_41461 = T_41460 & T_4334_82;
  assign T_41462 = T_41461 & T_4334_81;
  assign T_41463 = T_41462 & T_4334_80;
  assign T_41495 = T_41366 & T_4319_79;
  assign T_41527 = T_41398 & T_4324_79;
  assign T_41559 = T_41430 & T_4329_79;
  assign T_41591 = T_41462 & T_4334_79;
  assign T_41622 = T_41365 & T_4319_80;
  assign T_41623 = T_41622 & T_4319_79;
  assign T_41654 = T_41397 & T_4324_80;
  assign T_41655 = T_41654 & T_4324_79;
  assign T_41686 = T_41429 & T_4329_80;
  assign T_41687 = T_41686 & T_4329_79;
  assign T_41718 = T_41461 & T_4334_80;
  assign T_41719 = T_41718 & T_4334_79;
  assign T_41749 = T_41364 & T_4319_81;
  assign T_41750 = T_41749 & T_4319_80;
  assign T_41751 = T_41750 & T_4319_79;
  assign T_41781 = T_41396 & T_4324_81;
  assign T_41782 = T_41781 & T_4324_80;
  assign T_41783 = T_41782 & T_4324_79;
  assign T_41813 = T_41428 & T_4329_81;
  assign T_41814 = T_41813 & T_4329_80;
  assign T_41815 = T_41814 & T_4329_79;
  assign T_41845 = T_41460 & T_4334_81;
  assign T_41846 = T_41845 & T_4334_80;
  assign T_41847 = T_41846 & T_4334_79;
  assign T_41876 = T_41363 & T_4319_82;
  assign T_41877 = T_41876 & T_4319_81;
  assign T_41878 = T_41877 & T_4319_80;
  assign T_41879 = T_41878 & T_4319_79;
  assign T_41908 = T_41395 & T_4324_82;
  assign T_41909 = T_41908 & T_4324_81;
  assign T_41910 = T_41909 & T_4324_80;
  assign T_41911 = T_41910 & T_4324_79;
  assign T_41940 = T_41427 & T_4329_82;
  assign T_41941 = T_41940 & T_4329_81;
  assign T_41942 = T_41941 & T_4329_80;
  assign T_41943 = T_41942 & T_4329_79;
  assign T_41972 = T_41459 & T_4334_82;
  assign T_41973 = T_41972 & T_4334_81;
  assign T_41974 = T_41973 & T_4334_80;
  assign T_41975 = T_41974 & T_4334_79;
  assign T_42003 = T_41362 & T_4319_83;
  assign T_42004 = T_42003 & T_4319_82;
  assign T_42005 = T_42004 & T_4319_81;
  assign T_42006 = T_42005 & T_4319_80;
  assign T_42007 = T_42006 & T_4319_79;
  assign T_42035 = T_41394 & T_4324_83;
  assign T_42036 = T_42035 & T_4324_82;
  assign T_42037 = T_42036 & T_4324_81;
  assign T_42038 = T_42037 & T_4324_80;
  assign T_42039 = T_42038 & T_4324_79;
  assign T_42067 = T_41426 & T_4329_83;
  assign T_42068 = T_42067 & T_4329_82;
  assign T_42069 = T_42068 & T_4329_81;
  assign T_42070 = T_42069 & T_4329_80;
  assign T_42071 = T_42070 & T_4329_79;
  assign T_42099 = T_41458 & T_4334_83;
  assign T_42100 = T_42099 & T_4334_82;
  assign T_42101 = T_42100 & T_4334_81;
  assign T_42102 = T_42101 & T_4334_80;
  assign T_42103 = T_42102 & T_4334_79;
  assign T_42130 = T_41361 & T_4319_84;
  assign T_42131 = T_42130 & T_4319_83;
  assign T_42132 = T_42131 & T_4319_82;
  assign T_42133 = T_42132 & T_4319_81;
  assign T_42134 = T_42133 & T_4319_80;
  assign T_42135 = T_42134 & T_4319_79;
  assign T_42162 = T_41393 & T_4324_84;
  assign T_42163 = T_42162 & T_4324_83;
  assign T_42164 = T_42163 & T_4324_82;
  assign T_42165 = T_42164 & T_4324_81;
  assign T_42166 = T_42165 & T_4324_80;
  assign T_42167 = T_42166 & T_4324_79;
  assign T_42194 = T_41425 & T_4329_84;
  assign T_42195 = T_42194 & T_4329_83;
  assign T_42196 = T_42195 & T_4329_82;
  assign T_42197 = T_42196 & T_4329_81;
  assign T_42198 = T_42197 & T_4329_80;
  assign T_42199 = T_42198 & T_4329_79;
  assign T_42226 = T_41457 & T_4334_84;
  assign T_42227 = T_42226 & T_4334_83;
  assign T_42228 = T_42227 & T_4334_82;
  assign T_42229 = T_42228 & T_4334_81;
  assign T_42230 = T_42229 & T_4334_80;
  assign T_42231 = T_42230 & T_4334_79;
  assign T_42257 = T_41360 & T_4319_85;
  assign T_42258 = T_42257 & T_4319_84;
  assign T_42259 = T_42258 & T_4319_83;
  assign T_42260 = T_42259 & T_4319_82;
  assign T_42261 = T_42260 & T_4319_81;
  assign T_42262 = T_42261 & T_4319_80;
  assign T_42263 = T_42262 & T_4319_79;
  assign T_42289 = T_41392 & T_4324_85;
  assign T_42290 = T_42289 & T_4324_84;
  assign T_42291 = T_42290 & T_4324_83;
  assign T_42292 = T_42291 & T_4324_82;
  assign T_42293 = T_42292 & T_4324_81;
  assign T_42294 = T_42293 & T_4324_80;
  assign T_42295 = T_42294 & T_4324_79;
  assign T_42321 = T_41424 & T_4329_85;
  assign T_42322 = T_42321 & T_4329_84;
  assign T_42323 = T_42322 & T_4329_83;
  assign T_42324 = T_42323 & T_4329_82;
  assign T_42325 = T_42324 & T_4329_81;
  assign T_42326 = T_42325 & T_4329_80;
  assign T_42327 = T_42326 & T_4329_79;
  assign T_42353 = T_41456 & T_4334_85;
  assign T_42354 = T_42353 & T_4334_84;
  assign T_42355 = T_42354 & T_4334_83;
  assign T_42356 = T_42355 & T_4334_82;
  assign T_42357 = T_42356 & T_4334_81;
  assign T_42358 = T_42357 & T_4334_80;
  assign T_42359 = T_42358 & T_4334_79;
  assign T_42384 = T_41359 & T_4319_86;
  assign T_42385 = T_42384 & T_4319_85;
  assign T_42386 = T_42385 & T_4319_84;
  assign T_42387 = T_42386 & T_4319_83;
  assign T_42388 = T_42387 & T_4319_82;
  assign T_42389 = T_42388 & T_4319_81;
  assign T_42390 = T_42389 & T_4319_80;
  assign T_42391 = T_42390 & T_4319_79;
  assign T_42416 = T_41391 & T_4324_86;
  assign T_42417 = T_42416 & T_4324_85;
  assign T_42418 = T_42417 & T_4324_84;
  assign T_42419 = T_42418 & T_4324_83;
  assign T_42420 = T_42419 & T_4324_82;
  assign T_42421 = T_42420 & T_4324_81;
  assign T_42422 = T_42421 & T_4324_80;
  assign T_42423 = T_42422 & T_4324_79;
  assign T_42448 = T_41423 & T_4329_86;
  assign T_42449 = T_42448 & T_4329_85;
  assign T_42450 = T_42449 & T_4329_84;
  assign T_42451 = T_42450 & T_4329_83;
  assign T_42452 = T_42451 & T_4329_82;
  assign T_42453 = T_42452 & T_4329_81;
  assign T_42454 = T_42453 & T_4329_80;
  assign T_42455 = T_42454 & T_4329_79;
  assign T_42480 = T_41455 & T_4334_86;
  assign T_42481 = T_42480 & T_4334_85;
  assign T_42482 = T_42481 & T_4334_84;
  assign T_42483 = T_42482 & T_4334_83;
  assign T_42484 = T_42483 & T_4334_82;
  assign T_42485 = T_42484 & T_4334_81;
  assign T_42486 = T_42485 & T_4334_80;
  assign T_42487 = T_42486 & T_4334_79;
  assign T_42511 = T_41358 & T_4319_87;
  assign T_42512 = T_42511 & T_4319_86;
  assign T_42513 = T_42512 & T_4319_85;
  assign T_42514 = T_42513 & T_4319_84;
  assign T_42515 = T_42514 & T_4319_83;
  assign T_42516 = T_42515 & T_4319_82;
  assign T_42517 = T_42516 & T_4319_81;
  assign T_42518 = T_42517 & T_4319_80;
  assign T_42519 = T_42518 & T_4319_79;
  assign T_42543 = T_41390 & T_4324_87;
  assign T_42544 = T_42543 & T_4324_86;
  assign T_42545 = T_42544 & T_4324_85;
  assign T_42546 = T_42545 & T_4324_84;
  assign T_42547 = T_42546 & T_4324_83;
  assign T_42548 = T_42547 & T_4324_82;
  assign T_42549 = T_42548 & T_4324_81;
  assign T_42550 = T_42549 & T_4324_80;
  assign T_42551 = T_42550 & T_4324_79;
  assign T_42575 = T_41422 & T_4329_87;
  assign T_42576 = T_42575 & T_4329_86;
  assign T_42577 = T_42576 & T_4329_85;
  assign T_42578 = T_42577 & T_4329_84;
  assign T_42579 = T_42578 & T_4329_83;
  assign T_42580 = T_42579 & T_4329_82;
  assign T_42581 = T_42580 & T_4329_81;
  assign T_42582 = T_42581 & T_4329_80;
  assign T_42583 = T_42582 & T_4329_79;
  assign T_42607 = T_41454 & T_4334_87;
  assign T_42608 = T_42607 & T_4334_86;
  assign T_42609 = T_42608 & T_4334_85;
  assign T_42610 = T_42609 & T_4334_84;
  assign T_42611 = T_42610 & T_4334_83;
  assign T_42612 = T_42611 & T_4334_82;
  assign T_42613 = T_42612 & T_4334_81;
  assign T_42614 = T_42613 & T_4334_80;
  assign T_42615 = T_42614 & T_4334_79;
  assign T_42638 = T_41357 & T_4319_88;
  assign T_42639 = T_42638 & T_4319_87;
  assign T_42640 = T_42639 & T_4319_86;
  assign T_42641 = T_42640 & T_4319_85;
  assign T_42642 = T_42641 & T_4319_84;
  assign T_42643 = T_42642 & T_4319_83;
  assign T_42644 = T_42643 & T_4319_82;
  assign T_42645 = T_42644 & T_4319_81;
  assign T_42646 = T_42645 & T_4319_80;
  assign T_42647 = T_42646 & T_4319_79;
  assign T_42670 = T_41389 & T_4324_88;
  assign T_42671 = T_42670 & T_4324_87;
  assign T_42672 = T_42671 & T_4324_86;
  assign T_42673 = T_42672 & T_4324_85;
  assign T_42674 = T_42673 & T_4324_84;
  assign T_42675 = T_42674 & T_4324_83;
  assign T_42676 = T_42675 & T_4324_82;
  assign T_42677 = T_42676 & T_4324_81;
  assign T_42678 = T_42677 & T_4324_80;
  assign T_42679 = T_42678 & T_4324_79;
  assign T_42702 = T_41421 & T_4329_88;
  assign T_42703 = T_42702 & T_4329_87;
  assign T_42704 = T_42703 & T_4329_86;
  assign T_42705 = T_42704 & T_4329_85;
  assign T_42706 = T_42705 & T_4329_84;
  assign T_42707 = T_42706 & T_4329_83;
  assign T_42708 = T_42707 & T_4329_82;
  assign T_42709 = T_42708 & T_4329_81;
  assign T_42710 = T_42709 & T_4329_80;
  assign T_42711 = T_42710 & T_4329_79;
  assign T_42734 = T_41453 & T_4334_88;
  assign T_42735 = T_42734 & T_4334_87;
  assign T_42736 = T_42735 & T_4334_86;
  assign T_42737 = T_42736 & T_4334_85;
  assign T_42738 = T_42737 & T_4334_84;
  assign T_42739 = T_42738 & T_4334_83;
  assign T_42740 = T_42739 & T_4334_82;
  assign T_42741 = T_42740 & T_4334_81;
  assign T_42742 = T_42741 & T_4334_80;
  assign T_42743 = T_42742 & T_4334_79;
  assign T_42765 = T_41356 & T_4319_89;
  assign T_42766 = T_42765 & T_4319_88;
  assign T_42767 = T_42766 & T_4319_87;
  assign T_42768 = T_42767 & T_4319_86;
  assign T_42769 = T_42768 & T_4319_85;
  assign T_42770 = T_42769 & T_4319_84;
  assign T_42771 = T_42770 & T_4319_83;
  assign T_42772 = T_42771 & T_4319_82;
  assign T_42773 = T_42772 & T_4319_81;
  assign T_42774 = T_42773 & T_4319_80;
  assign T_42775 = T_42774 & T_4319_79;
  assign T_42797 = T_41388 & T_4324_89;
  assign T_42798 = T_42797 & T_4324_88;
  assign T_42799 = T_42798 & T_4324_87;
  assign T_42800 = T_42799 & T_4324_86;
  assign T_42801 = T_42800 & T_4324_85;
  assign T_42802 = T_42801 & T_4324_84;
  assign T_42803 = T_42802 & T_4324_83;
  assign T_42804 = T_42803 & T_4324_82;
  assign T_42805 = T_42804 & T_4324_81;
  assign T_42806 = T_42805 & T_4324_80;
  assign T_42807 = T_42806 & T_4324_79;
  assign T_42829 = T_41420 & T_4329_89;
  assign T_42830 = T_42829 & T_4329_88;
  assign T_42831 = T_42830 & T_4329_87;
  assign T_42832 = T_42831 & T_4329_86;
  assign T_42833 = T_42832 & T_4329_85;
  assign T_42834 = T_42833 & T_4329_84;
  assign T_42835 = T_42834 & T_4329_83;
  assign T_42836 = T_42835 & T_4329_82;
  assign T_42837 = T_42836 & T_4329_81;
  assign T_42838 = T_42837 & T_4329_80;
  assign T_42839 = T_42838 & T_4329_79;
  assign T_42861 = T_41452 & T_4334_89;
  assign T_42862 = T_42861 & T_4334_88;
  assign T_42863 = T_42862 & T_4334_87;
  assign T_42864 = T_42863 & T_4334_86;
  assign T_42865 = T_42864 & T_4334_85;
  assign T_42866 = T_42865 & T_4334_84;
  assign T_42867 = T_42866 & T_4334_83;
  assign T_42868 = T_42867 & T_4334_82;
  assign T_42869 = T_42868 & T_4334_81;
  assign T_42870 = T_42869 & T_4334_80;
  assign T_42871 = T_42870 & T_4334_79;
  assign T_42892 = T_41355 & T_4319_90;
  assign T_42893 = T_42892 & T_4319_89;
  assign T_42894 = T_42893 & T_4319_88;
  assign T_42895 = T_42894 & T_4319_87;
  assign T_42896 = T_42895 & T_4319_86;
  assign T_42897 = T_42896 & T_4319_85;
  assign T_42898 = T_42897 & T_4319_84;
  assign T_42899 = T_42898 & T_4319_83;
  assign T_42900 = T_42899 & T_4319_82;
  assign T_42901 = T_42900 & T_4319_81;
  assign T_42902 = T_42901 & T_4319_80;
  assign T_42903 = T_42902 & T_4319_79;
  assign T_42924 = T_41387 & T_4324_90;
  assign T_42925 = T_42924 & T_4324_89;
  assign T_42926 = T_42925 & T_4324_88;
  assign T_42927 = T_42926 & T_4324_87;
  assign T_42928 = T_42927 & T_4324_86;
  assign T_42929 = T_42928 & T_4324_85;
  assign T_42930 = T_42929 & T_4324_84;
  assign T_42931 = T_42930 & T_4324_83;
  assign T_42932 = T_42931 & T_4324_82;
  assign T_42933 = T_42932 & T_4324_81;
  assign T_42934 = T_42933 & T_4324_80;
  assign T_42935 = T_42934 & T_4324_79;
  assign T_42956 = T_41419 & T_4329_90;
  assign T_42957 = T_42956 & T_4329_89;
  assign T_42958 = T_42957 & T_4329_88;
  assign T_42959 = T_42958 & T_4329_87;
  assign T_42960 = T_42959 & T_4329_86;
  assign T_42961 = T_42960 & T_4329_85;
  assign T_42962 = T_42961 & T_4329_84;
  assign T_42963 = T_42962 & T_4329_83;
  assign T_42964 = T_42963 & T_4329_82;
  assign T_42965 = T_42964 & T_4329_81;
  assign T_42966 = T_42965 & T_4329_80;
  assign T_42967 = T_42966 & T_4329_79;
  assign T_42988 = T_41451 & T_4334_90;
  assign T_42989 = T_42988 & T_4334_89;
  assign T_42990 = T_42989 & T_4334_88;
  assign T_42991 = T_42990 & T_4334_87;
  assign T_42992 = T_42991 & T_4334_86;
  assign T_42993 = T_42992 & T_4334_85;
  assign T_42994 = T_42993 & T_4334_84;
  assign T_42995 = T_42994 & T_4334_83;
  assign T_42996 = T_42995 & T_4334_82;
  assign T_42997 = T_42996 & T_4334_81;
  assign T_42998 = T_42997 & T_4334_80;
  assign T_42999 = T_42998 & T_4334_79;
  assign T_43019 = T_41354 & T_4319_91;
  assign T_43020 = T_43019 & T_4319_90;
  assign T_43021 = T_43020 & T_4319_89;
  assign T_43022 = T_43021 & T_4319_88;
  assign T_43023 = T_43022 & T_4319_87;
  assign T_43024 = T_43023 & T_4319_86;
  assign T_43025 = T_43024 & T_4319_85;
  assign T_43026 = T_43025 & T_4319_84;
  assign T_43027 = T_43026 & T_4319_83;
  assign T_43028 = T_43027 & T_4319_82;
  assign T_43029 = T_43028 & T_4319_81;
  assign T_43030 = T_43029 & T_4319_80;
  assign T_43031 = T_43030 & T_4319_79;
  assign T_43051 = T_41386 & T_4324_91;
  assign T_43052 = T_43051 & T_4324_90;
  assign T_43053 = T_43052 & T_4324_89;
  assign T_43054 = T_43053 & T_4324_88;
  assign T_43055 = T_43054 & T_4324_87;
  assign T_43056 = T_43055 & T_4324_86;
  assign T_43057 = T_43056 & T_4324_85;
  assign T_43058 = T_43057 & T_4324_84;
  assign T_43059 = T_43058 & T_4324_83;
  assign T_43060 = T_43059 & T_4324_82;
  assign T_43061 = T_43060 & T_4324_81;
  assign T_43062 = T_43061 & T_4324_80;
  assign T_43063 = T_43062 & T_4324_79;
  assign T_43083 = T_41418 & T_4329_91;
  assign T_43084 = T_43083 & T_4329_90;
  assign T_43085 = T_43084 & T_4329_89;
  assign T_43086 = T_43085 & T_4329_88;
  assign T_43087 = T_43086 & T_4329_87;
  assign T_43088 = T_43087 & T_4329_86;
  assign T_43089 = T_43088 & T_4329_85;
  assign T_43090 = T_43089 & T_4329_84;
  assign T_43091 = T_43090 & T_4329_83;
  assign T_43092 = T_43091 & T_4329_82;
  assign T_43093 = T_43092 & T_4329_81;
  assign T_43094 = T_43093 & T_4329_80;
  assign T_43095 = T_43094 & T_4329_79;
  assign T_43115 = T_41450 & T_4334_91;
  assign T_43116 = T_43115 & T_4334_90;
  assign T_43117 = T_43116 & T_4334_89;
  assign T_43118 = T_43117 & T_4334_88;
  assign T_43119 = T_43118 & T_4334_87;
  assign T_43120 = T_43119 & T_4334_86;
  assign T_43121 = T_43120 & T_4334_85;
  assign T_43122 = T_43121 & T_4334_84;
  assign T_43123 = T_43122 & T_4334_83;
  assign T_43124 = T_43123 & T_4334_82;
  assign T_43125 = T_43124 & T_4334_81;
  assign T_43126 = T_43125 & T_4334_80;
  assign T_43127 = T_43126 & T_4334_79;
  assign T_43146 = T_41353 & T_4319_92;
  assign T_43147 = T_43146 & T_4319_91;
  assign T_43148 = T_43147 & T_4319_90;
  assign T_43149 = T_43148 & T_4319_89;
  assign T_43150 = T_43149 & T_4319_88;
  assign T_43151 = T_43150 & T_4319_87;
  assign T_43152 = T_43151 & T_4319_86;
  assign T_43153 = T_43152 & T_4319_85;
  assign T_43154 = T_43153 & T_4319_84;
  assign T_43155 = T_43154 & T_4319_83;
  assign T_43156 = T_43155 & T_4319_82;
  assign T_43157 = T_43156 & T_4319_81;
  assign T_43158 = T_43157 & T_4319_80;
  assign T_43159 = T_43158 & T_4319_79;
  assign T_43178 = T_41385 & T_4324_92;
  assign T_43179 = T_43178 & T_4324_91;
  assign T_43180 = T_43179 & T_4324_90;
  assign T_43181 = T_43180 & T_4324_89;
  assign T_43182 = T_43181 & T_4324_88;
  assign T_43183 = T_43182 & T_4324_87;
  assign T_43184 = T_43183 & T_4324_86;
  assign T_43185 = T_43184 & T_4324_85;
  assign T_43186 = T_43185 & T_4324_84;
  assign T_43187 = T_43186 & T_4324_83;
  assign T_43188 = T_43187 & T_4324_82;
  assign T_43189 = T_43188 & T_4324_81;
  assign T_43190 = T_43189 & T_4324_80;
  assign T_43191 = T_43190 & T_4324_79;
  assign T_43210 = T_41417 & T_4329_92;
  assign T_43211 = T_43210 & T_4329_91;
  assign T_43212 = T_43211 & T_4329_90;
  assign T_43213 = T_43212 & T_4329_89;
  assign T_43214 = T_43213 & T_4329_88;
  assign T_43215 = T_43214 & T_4329_87;
  assign T_43216 = T_43215 & T_4329_86;
  assign T_43217 = T_43216 & T_4329_85;
  assign T_43218 = T_43217 & T_4329_84;
  assign T_43219 = T_43218 & T_4329_83;
  assign T_43220 = T_43219 & T_4329_82;
  assign T_43221 = T_43220 & T_4329_81;
  assign T_43222 = T_43221 & T_4329_80;
  assign T_43223 = T_43222 & T_4329_79;
  assign T_43242 = T_41449 & T_4334_92;
  assign T_43243 = T_43242 & T_4334_91;
  assign T_43244 = T_43243 & T_4334_90;
  assign T_43245 = T_43244 & T_4334_89;
  assign T_43246 = T_43245 & T_4334_88;
  assign T_43247 = T_43246 & T_4334_87;
  assign T_43248 = T_43247 & T_4334_86;
  assign T_43249 = T_43248 & T_4334_85;
  assign T_43250 = T_43249 & T_4334_84;
  assign T_43251 = T_43250 & T_4334_83;
  assign T_43252 = T_43251 & T_4334_82;
  assign T_43253 = T_43252 & T_4334_81;
  assign T_43254 = T_43253 & T_4334_80;
  assign T_43255 = T_43254 & T_4334_79;
  assign T_43273 = T_41352 & T_4319_93;
  assign T_43274 = T_43273 & T_4319_92;
  assign T_43275 = T_43274 & T_4319_91;
  assign T_43276 = T_43275 & T_4319_90;
  assign T_43277 = T_43276 & T_4319_89;
  assign T_43278 = T_43277 & T_4319_88;
  assign T_43279 = T_43278 & T_4319_87;
  assign T_43280 = T_43279 & T_4319_86;
  assign T_43281 = T_43280 & T_4319_85;
  assign T_43282 = T_43281 & T_4319_84;
  assign T_43283 = T_43282 & T_4319_83;
  assign T_43284 = T_43283 & T_4319_82;
  assign T_43285 = T_43284 & T_4319_81;
  assign T_43286 = T_43285 & T_4319_80;
  assign T_43287 = T_43286 & T_4319_79;
  assign T_43305 = T_41384 & T_4324_93;
  assign T_43306 = T_43305 & T_4324_92;
  assign T_43307 = T_43306 & T_4324_91;
  assign T_43308 = T_43307 & T_4324_90;
  assign T_43309 = T_43308 & T_4324_89;
  assign T_43310 = T_43309 & T_4324_88;
  assign T_43311 = T_43310 & T_4324_87;
  assign T_43312 = T_43311 & T_4324_86;
  assign T_43313 = T_43312 & T_4324_85;
  assign T_43314 = T_43313 & T_4324_84;
  assign T_43315 = T_43314 & T_4324_83;
  assign T_43316 = T_43315 & T_4324_82;
  assign T_43317 = T_43316 & T_4324_81;
  assign T_43318 = T_43317 & T_4324_80;
  assign T_43319 = T_43318 & T_4324_79;
  assign T_43337 = T_41416 & T_4329_93;
  assign T_43338 = T_43337 & T_4329_92;
  assign T_43339 = T_43338 & T_4329_91;
  assign T_43340 = T_43339 & T_4329_90;
  assign T_43341 = T_43340 & T_4329_89;
  assign T_43342 = T_43341 & T_4329_88;
  assign T_43343 = T_43342 & T_4329_87;
  assign T_43344 = T_43343 & T_4329_86;
  assign T_43345 = T_43344 & T_4329_85;
  assign T_43346 = T_43345 & T_4329_84;
  assign T_43347 = T_43346 & T_4329_83;
  assign T_43348 = T_43347 & T_4329_82;
  assign T_43349 = T_43348 & T_4329_81;
  assign T_43350 = T_43349 & T_4329_80;
  assign T_43351 = T_43350 & T_4329_79;
  assign T_43369 = T_41448 & T_4334_93;
  assign T_43370 = T_43369 & T_4334_92;
  assign T_43371 = T_43370 & T_4334_91;
  assign T_43372 = T_43371 & T_4334_90;
  assign T_43373 = T_43372 & T_4334_89;
  assign T_43374 = T_43373 & T_4334_88;
  assign T_43375 = T_43374 & T_4334_87;
  assign T_43376 = T_43375 & T_4334_86;
  assign T_43377 = T_43376 & T_4334_85;
  assign T_43378 = T_43377 & T_4334_84;
  assign T_43379 = T_43378 & T_4334_83;
  assign T_43380 = T_43379 & T_4334_82;
  assign T_43381 = T_43380 & T_4334_81;
  assign T_43382 = T_43381 & T_4334_80;
  assign T_43383 = T_43382 & T_4334_79;
  assign T_43400 = T_41351 & T_4319_94;
  assign T_43401 = T_43400 & T_4319_93;
  assign T_43402 = T_43401 & T_4319_92;
  assign T_43403 = T_43402 & T_4319_91;
  assign T_43404 = T_43403 & T_4319_90;
  assign T_43405 = T_43404 & T_4319_89;
  assign T_43406 = T_43405 & T_4319_88;
  assign T_43407 = T_43406 & T_4319_87;
  assign T_43408 = T_43407 & T_4319_86;
  assign T_43409 = T_43408 & T_4319_85;
  assign T_43410 = T_43409 & T_4319_84;
  assign T_43411 = T_43410 & T_4319_83;
  assign T_43412 = T_43411 & T_4319_82;
  assign T_43413 = T_43412 & T_4319_81;
  assign T_43414 = T_43413 & T_4319_80;
  assign T_43415 = T_43414 & T_4319_79;
  assign T_43432 = T_41383 & T_4324_94;
  assign T_43433 = T_43432 & T_4324_93;
  assign T_43434 = T_43433 & T_4324_92;
  assign T_43435 = T_43434 & T_4324_91;
  assign T_43436 = T_43435 & T_4324_90;
  assign T_43437 = T_43436 & T_4324_89;
  assign T_43438 = T_43437 & T_4324_88;
  assign T_43439 = T_43438 & T_4324_87;
  assign T_43440 = T_43439 & T_4324_86;
  assign T_43441 = T_43440 & T_4324_85;
  assign T_43442 = T_43441 & T_4324_84;
  assign T_43443 = T_43442 & T_4324_83;
  assign T_43444 = T_43443 & T_4324_82;
  assign T_43445 = T_43444 & T_4324_81;
  assign T_43446 = T_43445 & T_4324_80;
  assign T_43447 = T_43446 & T_4324_79;
  assign T_43464 = T_41415 & T_4329_94;
  assign T_43465 = T_43464 & T_4329_93;
  assign T_43466 = T_43465 & T_4329_92;
  assign T_43467 = T_43466 & T_4329_91;
  assign T_43468 = T_43467 & T_4329_90;
  assign T_43469 = T_43468 & T_4329_89;
  assign T_43470 = T_43469 & T_4329_88;
  assign T_43471 = T_43470 & T_4329_87;
  assign T_43472 = T_43471 & T_4329_86;
  assign T_43473 = T_43472 & T_4329_85;
  assign T_43474 = T_43473 & T_4329_84;
  assign T_43475 = T_43474 & T_4329_83;
  assign T_43476 = T_43475 & T_4329_82;
  assign T_43477 = T_43476 & T_4329_81;
  assign T_43478 = T_43477 & T_4329_80;
  assign T_43479 = T_43478 & T_4329_79;
  assign T_43496 = T_41447 & T_4334_94;
  assign T_43497 = T_43496 & T_4334_93;
  assign T_43498 = T_43497 & T_4334_92;
  assign T_43499 = T_43498 & T_4334_91;
  assign T_43500 = T_43499 & T_4334_90;
  assign T_43501 = T_43500 & T_4334_89;
  assign T_43502 = T_43501 & T_4334_88;
  assign T_43503 = T_43502 & T_4334_87;
  assign T_43504 = T_43503 & T_4334_86;
  assign T_43505 = T_43504 & T_4334_85;
  assign T_43506 = T_43505 & T_4334_84;
  assign T_43507 = T_43506 & T_4334_83;
  assign T_43508 = T_43507 & T_4334_82;
  assign T_43509 = T_43508 & T_4334_81;
  assign T_43510 = T_43509 & T_4334_80;
  assign T_43511 = T_43510 & T_4334_79;
  assign T_43527 = T_41350 & T_4319_95;
  assign T_43528 = T_43527 & T_4319_94;
  assign T_43529 = T_43528 & T_4319_93;
  assign T_43530 = T_43529 & T_4319_92;
  assign T_43531 = T_43530 & T_4319_91;
  assign T_43532 = T_43531 & T_4319_90;
  assign T_43533 = T_43532 & T_4319_89;
  assign T_43534 = T_43533 & T_4319_88;
  assign T_43535 = T_43534 & T_4319_87;
  assign T_43536 = T_43535 & T_4319_86;
  assign T_43537 = T_43536 & T_4319_85;
  assign T_43538 = T_43537 & T_4319_84;
  assign T_43539 = T_43538 & T_4319_83;
  assign T_43540 = T_43539 & T_4319_82;
  assign T_43541 = T_43540 & T_4319_81;
  assign T_43542 = T_43541 & T_4319_80;
  assign T_43543 = T_43542 & T_4319_79;
  assign T_43559 = T_41382 & T_4324_95;
  assign T_43560 = T_43559 & T_4324_94;
  assign T_43561 = T_43560 & T_4324_93;
  assign T_43562 = T_43561 & T_4324_92;
  assign T_43563 = T_43562 & T_4324_91;
  assign T_43564 = T_43563 & T_4324_90;
  assign T_43565 = T_43564 & T_4324_89;
  assign T_43566 = T_43565 & T_4324_88;
  assign T_43567 = T_43566 & T_4324_87;
  assign T_43568 = T_43567 & T_4324_86;
  assign T_43569 = T_43568 & T_4324_85;
  assign T_43570 = T_43569 & T_4324_84;
  assign T_43571 = T_43570 & T_4324_83;
  assign T_43572 = T_43571 & T_4324_82;
  assign T_43573 = T_43572 & T_4324_81;
  assign T_43574 = T_43573 & T_4324_80;
  assign T_43575 = T_43574 & T_4324_79;
  assign T_43591 = T_41414 & T_4329_95;
  assign T_43592 = T_43591 & T_4329_94;
  assign T_43593 = T_43592 & T_4329_93;
  assign T_43594 = T_43593 & T_4329_92;
  assign T_43595 = T_43594 & T_4329_91;
  assign T_43596 = T_43595 & T_4329_90;
  assign T_43597 = T_43596 & T_4329_89;
  assign T_43598 = T_43597 & T_4329_88;
  assign T_43599 = T_43598 & T_4329_87;
  assign T_43600 = T_43599 & T_4329_86;
  assign T_43601 = T_43600 & T_4329_85;
  assign T_43602 = T_43601 & T_4329_84;
  assign T_43603 = T_43602 & T_4329_83;
  assign T_43604 = T_43603 & T_4329_82;
  assign T_43605 = T_43604 & T_4329_81;
  assign T_43606 = T_43605 & T_4329_80;
  assign T_43607 = T_43606 & T_4329_79;
  assign T_43623 = T_41446 & T_4334_95;
  assign T_43624 = T_43623 & T_4334_94;
  assign T_43625 = T_43624 & T_4334_93;
  assign T_43626 = T_43625 & T_4334_92;
  assign T_43627 = T_43626 & T_4334_91;
  assign T_43628 = T_43627 & T_4334_90;
  assign T_43629 = T_43628 & T_4334_89;
  assign T_43630 = T_43629 & T_4334_88;
  assign T_43631 = T_43630 & T_4334_87;
  assign T_43632 = T_43631 & T_4334_86;
  assign T_43633 = T_43632 & T_4334_85;
  assign T_43634 = T_43633 & T_4334_84;
  assign T_43635 = T_43634 & T_4334_83;
  assign T_43636 = T_43635 & T_4334_82;
  assign T_43637 = T_43636 & T_4334_81;
  assign T_43638 = T_43637 & T_4334_80;
  assign T_43639 = T_43638 & T_4334_79;
  assign T_43654 = T_41349 & T_4319_96;
  assign T_43655 = T_43654 & T_4319_95;
  assign T_43656 = T_43655 & T_4319_94;
  assign T_43657 = T_43656 & T_4319_93;
  assign T_43658 = T_43657 & T_4319_92;
  assign T_43659 = T_43658 & T_4319_91;
  assign T_43660 = T_43659 & T_4319_90;
  assign T_43661 = T_43660 & T_4319_89;
  assign T_43662 = T_43661 & T_4319_88;
  assign T_43663 = T_43662 & T_4319_87;
  assign T_43664 = T_43663 & T_4319_86;
  assign T_43665 = T_43664 & T_4319_85;
  assign T_43666 = T_43665 & T_4319_84;
  assign T_43667 = T_43666 & T_4319_83;
  assign T_43668 = T_43667 & T_4319_82;
  assign T_43669 = T_43668 & T_4319_81;
  assign T_43670 = T_43669 & T_4319_80;
  assign T_43671 = T_43670 & T_4319_79;
  assign T_43686 = T_41381 & T_4324_96;
  assign T_43687 = T_43686 & T_4324_95;
  assign T_43688 = T_43687 & T_4324_94;
  assign T_43689 = T_43688 & T_4324_93;
  assign T_43690 = T_43689 & T_4324_92;
  assign T_43691 = T_43690 & T_4324_91;
  assign T_43692 = T_43691 & T_4324_90;
  assign T_43693 = T_43692 & T_4324_89;
  assign T_43694 = T_43693 & T_4324_88;
  assign T_43695 = T_43694 & T_4324_87;
  assign T_43696 = T_43695 & T_4324_86;
  assign T_43697 = T_43696 & T_4324_85;
  assign T_43698 = T_43697 & T_4324_84;
  assign T_43699 = T_43698 & T_4324_83;
  assign T_43700 = T_43699 & T_4324_82;
  assign T_43701 = T_43700 & T_4324_81;
  assign T_43702 = T_43701 & T_4324_80;
  assign T_43703 = T_43702 & T_4324_79;
  assign T_43718 = T_41413 & T_4329_96;
  assign T_43719 = T_43718 & T_4329_95;
  assign T_43720 = T_43719 & T_4329_94;
  assign T_43721 = T_43720 & T_4329_93;
  assign T_43722 = T_43721 & T_4329_92;
  assign T_43723 = T_43722 & T_4329_91;
  assign T_43724 = T_43723 & T_4329_90;
  assign T_43725 = T_43724 & T_4329_89;
  assign T_43726 = T_43725 & T_4329_88;
  assign T_43727 = T_43726 & T_4329_87;
  assign T_43728 = T_43727 & T_4329_86;
  assign T_43729 = T_43728 & T_4329_85;
  assign T_43730 = T_43729 & T_4329_84;
  assign T_43731 = T_43730 & T_4329_83;
  assign T_43732 = T_43731 & T_4329_82;
  assign T_43733 = T_43732 & T_4329_81;
  assign T_43734 = T_43733 & T_4329_80;
  assign T_43735 = T_43734 & T_4329_79;
  assign T_43750 = T_41445 & T_4334_96;
  assign T_43751 = T_43750 & T_4334_95;
  assign T_43752 = T_43751 & T_4334_94;
  assign T_43753 = T_43752 & T_4334_93;
  assign T_43754 = T_43753 & T_4334_92;
  assign T_43755 = T_43754 & T_4334_91;
  assign T_43756 = T_43755 & T_4334_90;
  assign T_43757 = T_43756 & T_4334_89;
  assign T_43758 = T_43757 & T_4334_88;
  assign T_43759 = T_43758 & T_4334_87;
  assign T_43760 = T_43759 & T_4334_86;
  assign T_43761 = T_43760 & T_4334_85;
  assign T_43762 = T_43761 & T_4334_84;
  assign T_43763 = T_43762 & T_4334_83;
  assign T_43764 = T_43763 & T_4334_82;
  assign T_43765 = T_43764 & T_4334_81;
  assign T_43766 = T_43765 & T_4334_80;
  assign T_43767 = T_43766 & T_4334_79;
  assign T_43781 = T_41348 & T_4319_97;
  assign T_43782 = T_43781 & T_4319_96;
  assign T_43783 = T_43782 & T_4319_95;
  assign T_43784 = T_43783 & T_4319_94;
  assign T_43785 = T_43784 & T_4319_93;
  assign T_43786 = T_43785 & T_4319_92;
  assign T_43787 = T_43786 & T_4319_91;
  assign T_43788 = T_43787 & T_4319_90;
  assign T_43789 = T_43788 & T_4319_89;
  assign T_43790 = T_43789 & T_4319_88;
  assign T_43791 = T_43790 & T_4319_87;
  assign T_43792 = T_43791 & T_4319_86;
  assign T_43793 = T_43792 & T_4319_85;
  assign T_43794 = T_43793 & T_4319_84;
  assign T_43795 = T_43794 & T_4319_83;
  assign T_43796 = T_43795 & T_4319_82;
  assign T_43797 = T_43796 & T_4319_81;
  assign T_43798 = T_43797 & T_4319_80;
  assign T_43799 = T_43798 & T_4319_79;
  assign T_43813 = T_41380 & T_4324_97;
  assign T_43814 = T_43813 & T_4324_96;
  assign T_43815 = T_43814 & T_4324_95;
  assign T_43816 = T_43815 & T_4324_94;
  assign T_43817 = T_43816 & T_4324_93;
  assign T_43818 = T_43817 & T_4324_92;
  assign T_43819 = T_43818 & T_4324_91;
  assign T_43820 = T_43819 & T_4324_90;
  assign T_43821 = T_43820 & T_4324_89;
  assign T_43822 = T_43821 & T_4324_88;
  assign T_43823 = T_43822 & T_4324_87;
  assign T_43824 = T_43823 & T_4324_86;
  assign T_43825 = T_43824 & T_4324_85;
  assign T_43826 = T_43825 & T_4324_84;
  assign T_43827 = T_43826 & T_4324_83;
  assign T_43828 = T_43827 & T_4324_82;
  assign T_43829 = T_43828 & T_4324_81;
  assign T_43830 = T_43829 & T_4324_80;
  assign T_43831 = T_43830 & T_4324_79;
  assign T_43845 = T_41412 & T_4329_97;
  assign T_43846 = T_43845 & T_4329_96;
  assign T_43847 = T_43846 & T_4329_95;
  assign T_43848 = T_43847 & T_4329_94;
  assign T_43849 = T_43848 & T_4329_93;
  assign T_43850 = T_43849 & T_4329_92;
  assign T_43851 = T_43850 & T_4329_91;
  assign T_43852 = T_43851 & T_4329_90;
  assign T_43853 = T_43852 & T_4329_89;
  assign T_43854 = T_43853 & T_4329_88;
  assign T_43855 = T_43854 & T_4329_87;
  assign T_43856 = T_43855 & T_4329_86;
  assign T_43857 = T_43856 & T_4329_85;
  assign T_43858 = T_43857 & T_4329_84;
  assign T_43859 = T_43858 & T_4329_83;
  assign T_43860 = T_43859 & T_4329_82;
  assign T_43861 = T_43860 & T_4329_81;
  assign T_43862 = T_43861 & T_4329_80;
  assign T_43863 = T_43862 & T_4329_79;
  assign T_43877 = T_41444 & T_4334_97;
  assign T_43878 = T_43877 & T_4334_96;
  assign T_43879 = T_43878 & T_4334_95;
  assign T_43880 = T_43879 & T_4334_94;
  assign T_43881 = T_43880 & T_4334_93;
  assign T_43882 = T_43881 & T_4334_92;
  assign T_43883 = T_43882 & T_4334_91;
  assign T_43884 = T_43883 & T_4334_90;
  assign T_43885 = T_43884 & T_4334_89;
  assign T_43886 = T_43885 & T_4334_88;
  assign T_43887 = T_43886 & T_4334_87;
  assign T_43888 = T_43887 & T_4334_86;
  assign T_43889 = T_43888 & T_4334_85;
  assign T_43890 = T_43889 & T_4334_84;
  assign T_43891 = T_43890 & T_4334_83;
  assign T_43892 = T_43891 & T_4334_82;
  assign T_43893 = T_43892 & T_4334_81;
  assign T_43894 = T_43893 & T_4334_80;
  assign T_43895 = T_43894 & T_4334_79;
  assign T_43908 = T_41347 & T_4319_98;
  assign T_43909 = T_43908 & T_4319_97;
  assign T_43910 = T_43909 & T_4319_96;
  assign T_43911 = T_43910 & T_4319_95;
  assign T_43912 = T_43911 & T_4319_94;
  assign T_43913 = T_43912 & T_4319_93;
  assign T_43914 = T_43913 & T_4319_92;
  assign T_43915 = T_43914 & T_4319_91;
  assign T_43916 = T_43915 & T_4319_90;
  assign T_43917 = T_43916 & T_4319_89;
  assign T_43918 = T_43917 & T_4319_88;
  assign T_43919 = T_43918 & T_4319_87;
  assign T_43920 = T_43919 & T_4319_86;
  assign T_43921 = T_43920 & T_4319_85;
  assign T_43922 = T_43921 & T_4319_84;
  assign T_43923 = T_43922 & T_4319_83;
  assign T_43924 = T_43923 & T_4319_82;
  assign T_43925 = T_43924 & T_4319_81;
  assign T_43926 = T_43925 & T_4319_80;
  assign T_43927 = T_43926 & T_4319_79;
  assign T_43940 = T_41379 & T_4324_98;
  assign T_43941 = T_43940 & T_4324_97;
  assign T_43942 = T_43941 & T_4324_96;
  assign T_43943 = T_43942 & T_4324_95;
  assign T_43944 = T_43943 & T_4324_94;
  assign T_43945 = T_43944 & T_4324_93;
  assign T_43946 = T_43945 & T_4324_92;
  assign T_43947 = T_43946 & T_4324_91;
  assign T_43948 = T_43947 & T_4324_90;
  assign T_43949 = T_43948 & T_4324_89;
  assign T_43950 = T_43949 & T_4324_88;
  assign T_43951 = T_43950 & T_4324_87;
  assign T_43952 = T_43951 & T_4324_86;
  assign T_43953 = T_43952 & T_4324_85;
  assign T_43954 = T_43953 & T_4324_84;
  assign T_43955 = T_43954 & T_4324_83;
  assign T_43956 = T_43955 & T_4324_82;
  assign T_43957 = T_43956 & T_4324_81;
  assign T_43958 = T_43957 & T_4324_80;
  assign T_43959 = T_43958 & T_4324_79;
  assign T_43972 = T_41411 & T_4329_98;
  assign T_43973 = T_43972 & T_4329_97;
  assign T_43974 = T_43973 & T_4329_96;
  assign T_43975 = T_43974 & T_4329_95;
  assign T_43976 = T_43975 & T_4329_94;
  assign T_43977 = T_43976 & T_4329_93;
  assign T_43978 = T_43977 & T_4329_92;
  assign T_43979 = T_43978 & T_4329_91;
  assign T_43980 = T_43979 & T_4329_90;
  assign T_43981 = T_43980 & T_4329_89;
  assign T_43982 = T_43981 & T_4329_88;
  assign T_43983 = T_43982 & T_4329_87;
  assign T_43984 = T_43983 & T_4329_86;
  assign T_43985 = T_43984 & T_4329_85;
  assign T_43986 = T_43985 & T_4329_84;
  assign T_43987 = T_43986 & T_4329_83;
  assign T_43988 = T_43987 & T_4329_82;
  assign T_43989 = T_43988 & T_4329_81;
  assign T_43990 = T_43989 & T_4329_80;
  assign T_43991 = T_43990 & T_4329_79;
  assign T_44004 = T_41443 & T_4334_98;
  assign T_44005 = T_44004 & T_4334_97;
  assign T_44006 = T_44005 & T_4334_96;
  assign T_44007 = T_44006 & T_4334_95;
  assign T_44008 = T_44007 & T_4334_94;
  assign T_44009 = T_44008 & T_4334_93;
  assign T_44010 = T_44009 & T_4334_92;
  assign T_44011 = T_44010 & T_4334_91;
  assign T_44012 = T_44011 & T_4334_90;
  assign T_44013 = T_44012 & T_4334_89;
  assign T_44014 = T_44013 & T_4334_88;
  assign T_44015 = T_44014 & T_4334_87;
  assign T_44016 = T_44015 & T_4334_86;
  assign T_44017 = T_44016 & T_4334_85;
  assign T_44018 = T_44017 & T_4334_84;
  assign T_44019 = T_44018 & T_4334_83;
  assign T_44020 = T_44019 & T_4334_82;
  assign T_44021 = T_44020 & T_4334_81;
  assign T_44022 = T_44021 & T_4334_80;
  assign T_44023 = T_44022 & T_4334_79;
  assign T_44035 = T_41346 & T_4319_99;
  assign T_44036 = T_44035 & T_4319_98;
  assign T_44037 = T_44036 & T_4319_97;
  assign T_44038 = T_44037 & T_4319_96;
  assign T_44039 = T_44038 & T_4319_95;
  assign T_44040 = T_44039 & T_4319_94;
  assign T_44041 = T_44040 & T_4319_93;
  assign T_44042 = T_44041 & T_4319_92;
  assign T_44043 = T_44042 & T_4319_91;
  assign T_44044 = T_44043 & T_4319_90;
  assign T_44045 = T_44044 & T_4319_89;
  assign T_44046 = T_44045 & T_4319_88;
  assign T_44047 = T_44046 & T_4319_87;
  assign T_44048 = T_44047 & T_4319_86;
  assign T_44049 = T_44048 & T_4319_85;
  assign T_44050 = T_44049 & T_4319_84;
  assign T_44051 = T_44050 & T_4319_83;
  assign T_44052 = T_44051 & T_4319_82;
  assign T_44053 = T_44052 & T_4319_81;
  assign T_44054 = T_44053 & T_4319_80;
  assign T_44055 = T_44054 & T_4319_79;
  assign T_44067 = T_41378 & T_4324_99;
  assign T_44068 = T_44067 & T_4324_98;
  assign T_44069 = T_44068 & T_4324_97;
  assign T_44070 = T_44069 & T_4324_96;
  assign T_44071 = T_44070 & T_4324_95;
  assign T_44072 = T_44071 & T_4324_94;
  assign T_44073 = T_44072 & T_4324_93;
  assign T_44074 = T_44073 & T_4324_92;
  assign T_44075 = T_44074 & T_4324_91;
  assign T_44076 = T_44075 & T_4324_90;
  assign T_44077 = T_44076 & T_4324_89;
  assign T_44078 = T_44077 & T_4324_88;
  assign T_44079 = T_44078 & T_4324_87;
  assign T_44080 = T_44079 & T_4324_86;
  assign T_44081 = T_44080 & T_4324_85;
  assign T_44082 = T_44081 & T_4324_84;
  assign T_44083 = T_44082 & T_4324_83;
  assign T_44084 = T_44083 & T_4324_82;
  assign T_44085 = T_44084 & T_4324_81;
  assign T_44086 = T_44085 & T_4324_80;
  assign T_44087 = T_44086 & T_4324_79;
  assign T_44099 = T_41410 & T_4329_99;
  assign T_44100 = T_44099 & T_4329_98;
  assign T_44101 = T_44100 & T_4329_97;
  assign T_44102 = T_44101 & T_4329_96;
  assign T_44103 = T_44102 & T_4329_95;
  assign T_44104 = T_44103 & T_4329_94;
  assign T_44105 = T_44104 & T_4329_93;
  assign T_44106 = T_44105 & T_4329_92;
  assign T_44107 = T_44106 & T_4329_91;
  assign T_44108 = T_44107 & T_4329_90;
  assign T_44109 = T_44108 & T_4329_89;
  assign T_44110 = T_44109 & T_4329_88;
  assign T_44111 = T_44110 & T_4329_87;
  assign T_44112 = T_44111 & T_4329_86;
  assign T_44113 = T_44112 & T_4329_85;
  assign T_44114 = T_44113 & T_4329_84;
  assign T_44115 = T_44114 & T_4329_83;
  assign T_44116 = T_44115 & T_4329_82;
  assign T_44117 = T_44116 & T_4329_81;
  assign T_44118 = T_44117 & T_4329_80;
  assign T_44119 = T_44118 & T_4329_79;
  assign T_44131 = T_41442 & T_4334_99;
  assign T_44132 = T_44131 & T_4334_98;
  assign T_44133 = T_44132 & T_4334_97;
  assign T_44134 = T_44133 & T_4334_96;
  assign T_44135 = T_44134 & T_4334_95;
  assign T_44136 = T_44135 & T_4334_94;
  assign T_44137 = T_44136 & T_4334_93;
  assign T_44138 = T_44137 & T_4334_92;
  assign T_44139 = T_44138 & T_4334_91;
  assign T_44140 = T_44139 & T_4334_90;
  assign T_44141 = T_44140 & T_4334_89;
  assign T_44142 = T_44141 & T_4334_88;
  assign T_44143 = T_44142 & T_4334_87;
  assign T_44144 = T_44143 & T_4334_86;
  assign T_44145 = T_44144 & T_4334_85;
  assign T_44146 = T_44145 & T_4334_84;
  assign T_44147 = T_44146 & T_4334_83;
  assign T_44148 = T_44147 & T_4334_82;
  assign T_44149 = T_44148 & T_4334_81;
  assign T_44150 = T_44149 & T_4334_80;
  assign T_44151 = T_44150 & T_4334_79;
  assign T_44162 = T_41345 & T_4319_100;
  assign T_44163 = T_44162 & T_4319_99;
  assign T_44164 = T_44163 & T_4319_98;
  assign T_44165 = T_44164 & T_4319_97;
  assign T_44166 = T_44165 & T_4319_96;
  assign T_44167 = T_44166 & T_4319_95;
  assign T_44168 = T_44167 & T_4319_94;
  assign T_44169 = T_44168 & T_4319_93;
  assign T_44170 = T_44169 & T_4319_92;
  assign T_44171 = T_44170 & T_4319_91;
  assign T_44172 = T_44171 & T_4319_90;
  assign T_44173 = T_44172 & T_4319_89;
  assign T_44174 = T_44173 & T_4319_88;
  assign T_44175 = T_44174 & T_4319_87;
  assign T_44176 = T_44175 & T_4319_86;
  assign T_44177 = T_44176 & T_4319_85;
  assign T_44178 = T_44177 & T_4319_84;
  assign T_44179 = T_44178 & T_4319_83;
  assign T_44180 = T_44179 & T_4319_82;
  assign T_44181 = T_44180 & T_4319_81;
  assign T_44182 = T_44181 & T_4319_80;
  assign T_44183 = T_44182 & T_4319_79;
  assign T_44194 = T_41377 & T_4324_100;
  assign T_44195 = T_44194 & T_4324_99;
  assign T_44196 = T_44195 & T_4324_98;
  assign T_44197 = T_44196 & T_4324_97;
  assign T_44198 = T_44197 & T_4324_96;
  assign T_44199 = T_44198 & T_4324_95;
  assign T_44200 = T_44199 & T_4324_94;
  assign T_44201 = T_44200 & T_4324_93;
  assign T_44202 = T_44201 & T_4324_92;
  assign T_44203 = T_44202 & T_4324_91;
  assign T_44204 = T_44203 & T_4324_90;
  assign T_44205 = T_44204 & T_4324_89;
  assign T_44206 = T_44205 & T_4324_88;
  assign T_44207 = T_44206 & T_4324_87;
  assign T_44208 = T_44207 & T_4324_86;
  assign T_44209 = T_44208 & T_4324_85;
  assign T_44210 = T_44209 & T_4324_84;
  assign T_44211 = T_44210 & T_4324_83;
  assign T_44212 = T_44211 & T_4324_82;
  assign T_44213 = T_44212 & T_4324_81;
  assign T_44214 = T_44213 & T_4324_80;
  assign T_44215 = T_44214 & T_4324_79;
  assign T_44226 = T_41409 & T_4329_100;
  assign T_44227 = T_44226 & T_4329_99;
  assign T_44228 = T_44227 & T_4329_98;
  assign T_44229 = T_44228 & T_4329_97;
  assign T_44230 = T_44229 & T_4329_96;
  assign T_44231 = T_44230 & T_4329_95;
  assign T_44232 = T_44231 & T_4329_94;
  assign T_44233 = T_44232 & T_4329_93;
  assign T_44234 = T_44233 & T_4329_92;
  assign T_44235 = T_44234 & T_4329_91;
  assign T_44236 = T_44235 & T_4329_90;
  assign T_44237 = T_44236 & T_4329_89;
  assign T_44238 = T_44237 & T_4329_88;
  assign T_44239 = T_44238 & T_4329_87;
  assign T_44240 = T_44239 & T_4329_86;
  assign T_44241 = T_44240 & T_4329_85;
  assign T_44242 = T_44241 & T_4329_84;
  assign T_44243 = T_44242 & T_4329_83;
  assign T_44244 = T_44243 & T_4329_82;
  assign T_44245 = T_44244 & T_4329_81;
  assign T_44246 = T_44245 & T_4329_80;
  assign T_44247 = T_44246 & T_4329_79;
  assign T_44258 = T_41441 & T_4334_100;
  assign T_44259 = T_44258 & T_4334_99;
  assign T_44260 = T_44259 & T_4334_98;
  assign T_44261 = T_44260 & T_4334_97;
  assign T_44262 = T_44261 & T_4334_96;
  assign T_44263 = T_44262 & T_4334_95;
  assign T_44264 = T_44263 & T_4334_94;
  assign T_44265 = T_44264 & T_4334_93;
  assign T_44266 = T_44265 & T_4334_92;
  assign T_44267 = T_44266 & T_4334_91;
  assign T_44268 = T_44267 & T_4334_90;
  assign T_44269 = T_44268 & T_4334_89;
  assign T_44270 = T_44269 & T_4334_88;
  assign T_44271 = T_44270 & T_4334_87;
  assign T_44272 = T_44271 & T_4334_86;
  assign T_44273 = T_44272 & T_4334_85;
  assign T_44274 = T_44273 & T_4334_84;
  assign T_44275 = T_44274 & T_4334_83;
  assign T_44276 = T_44275 & T_4334_82;
  assign T_44277 = T_44276 & T_4334_81;
  assign T_44278 = T_44277 & T_4334_80;
  assign T_44279 = T_44278 & T_4334_79;
  assign T_44289 = T_41344 & T_4319_101;
  assign T_44290 = T_44289 & T_4319_100;
  assign T_44291 = T_44290 & T_4319_99;
  assign T_44292 = T_44291 & T_4319_98;
  assign T_44293 = T_44292 & T_4319_97;
  assign T_44294 = T_44293 & T_4319_96;
  assign T_44295 = T_44294 & T_4319_95;
  assign T_44296 = T_44295 & T_4319_94;
  assign T_44297 = T_44296 & T_4319_93;
  assign T_44298 = T_44297 & T_4319_92;
  assign T_44299 = T_44298 & T_4319_91;
  assign T_44300 = T_44299 & T_4319_90;
  assign T_44301 = T_44300 & T_4319_89;
  assign T_44302 = T_44301 & T_4319_88;
  assign T_44303 = T_44302 & T_4319_87;
  assign T_44304 = T_44303 & T_4319_86;
  assign T_44305 = T_44304 & T_4319_85;
  assign T_44306 = T_44305 & T_4319_84;
  assign T_44307 = T_44306 & T_4319_83;
  assign T_44308 = T_44307 & T_4319_82;
  assign T_44309 = T_44308 & T_4319_81;
  assign T_44310 = T_44309 & T_4319_80;
  assign T_44311 = T_44310 & T_4319_79;
  assign T_44321 = T_41376 & T_4324_101;
  assign T_44322 = T_44321 & T_4324_100;
  assign T_44323 = T_44322 & T_4324_99;
  assign T_44324 = T_44323 & T_4324_98;
  assign T_44325 = T_44324 & T_4324_97;
  assign T_44326 = T_44325 & T_4324_96;
  assign T_44327 = T_44326 & T_4324_95;
  assign T_44328 = T_44327 & T_4324_94;
  assign T_44329 = T_44328 & T_4324_93;
  assign T_44330 = T_44329 & T_4324_92;
  assign T_44331 = T_44330 & T_4324_91;
  assign T_44332 = T_44331 & T_4324_90;
  assign T_44333 = T_44332 & T_4324_89;
  assign T_44334 = T_44333 & T_4324_88;
  assign T_44335 = T_44334 & T_4324_87;
  assign T_44336 = T_44335 & T_4324_86;
  assign T_44337 = T_44336 & T_4324_85;
  assign T_44338 = T_44337 & T_4324_84;
  assign T_44339 = T_44338 & T_4324_83;
  assign T_44340 = T_44339 & T_4324_82;
  assign T_44341 = T_44340 & T_4324_81;
  assign T_44342 = T_44341 & T_4324_80;
  assign T_44343 = T_44342 & T_4324_79;
  assign T_44353 = T_41408 & T_4329_101;
  assign T_44354 = T_44353 & T_4329_100;
  assign T_44355 = T_44354 & T_4329_99;
  assign T_44356 = T_44355 & T_4329_98;
  assign T_44357 = T_44356 & T_4329_97;
  assign T_44358 = T_44357 & T_4329_96;
  assign T_44359 = T_44358 & T_4329_95;
  assign T_44360 = T_44359 & T_4329_94;
  assign T_44361 = T_44360 & T_4329_93;
  assign T_44362 = T_44361 & T_4329_92;
  assign T_44363 = T_44362 & T_4329_91;
  assign T_44364 = T_44363 & T_4329_90;
  assign T_44365 = T_44364 & T_4329_89;
  assign T_44366 = T_44365 & T_4329_88;
  assign T_44367 = T_44366 & T_4329_87;
  assign T_44368 = T_44367 & T_4329_86;
  assign T_44369 = T_44368 & T_4329_85;
  assign T_44370 = T_44369 & T_4329_84;
  assign T_44371 = T_44370 & T_4329_83;
  assign T_44372 = T_44371 & T_4329_82;
  assign T_44373 = T_44372 & T_4329_81;
  assign T_44374 = T_44373 & T_4329_80;
  assign T_44375 = T_44374 & T_4329_79;
  assign T_44385 = T_41440 & T_4334_101;
  assign T_44386 = T_44385 & T_4334_100;
  assign T_44387 = T_44386 & T_4334_99;
  assign T_44388 = T_44387 & T_4334_98;
  assign T_44389 = T_44388 & T_4334_97;
  assign T_44390 = T_44389 & T_4334_96;
  assign T_44391 = T_44390 & T_4334_95;
  assign T_44392 = T_44391 & T_4334_94;
  assign T_44393 = T_44392 & T_4334_93;
  assign T_44394 = T_44393 & T_4334_92;
  assign T_44395 = T_44394 & T_4334_91;
  assign T_44396 = T_44395 & T_4334_90;
  assign T_44397 = T_44396 & T_4334_89;
  assign T_44398 = T_44397 & T_4334_88;
  assign T_44399 = T_44398 & T_4334_87;
  assign T_44400 = T_44399 & T_4334_86;
  assign T_44401 = T_44400 & T_4334_85;
  assign T_44402 = T_44401 & T_4334_84;
  assign T_44403 = T_44402 & T_4334_83;
  assign T_44404 = T_44403 & T_4334_82;
  assign T_44405 = T_44404 & T_4334_81;
  assign T_44406 = T_44405 & T_4334_80;
  assign T_44407 = T_44406 & T_4334_79;
  assign T_44416 = T_41343 & T_4319_102;
  assign T_44417 = T_44416 & T_4319_101;
  assign T_44418 = T_44417 & T_4319_100;
  assign T_44419 = T_44418 & T_4319_99;
  assign T_44420 = T_44419 & T_4319_98;
  assign T_44421 = T_44420 & T_4319_97;
  assign T_44422 = T_44421 & T_4319_96;
  assign T_44423 = T_44422 & T_4319_95;
  assign T_44424 = T_44423 & T_4319_94;
  assign T_44425 = T_44424 & T_4319_93;
  assign T_44426 = T_44425 & T_4319_92;
  assign T_44427 = T_44426 & T_4319_91;
  assign T_44428 = T_44427 & T_4319_90;
  assign T_44429 = T_44428 & T_4319_89;
  assign T_44430 = T_44429 & T_4319_88;
  assign T_44431 = T_44430 & T_4319_87;
  assign T_44432 = T_44431 & T_4319_86;
  assign T_44433 = T_44432 & T_4319_85;
  assign T_44434 = T_44433 & T_4319_84;
  assign T_44435 = T_44434 & T_4319_83;
  assign T_44436 = T_44435 & T_4319_82;
  assign T_44437 = T_44436 & T_4319_81;
  assign T_44438 = T_44437 & T_4319_80;
  assign T_44439 = T_44438 & T_4319_79;
  assign T_44448 = T_41375 & T_4324_102;
  assign T_44449 = T_44448 & T_4324_101;
  assign T_44450 = T_44449 & T_4324_100;
  assign T_44451 = T_44450 & T_4324_99;
  assign T_44452 = T_44451 & T_4324_98;
  assign T_44453 = T_44452 & T_4324_97;
  assign T_44454 = T_44453 & T_4324_96;
  assign T_44455 = T_44454 & T_4324_95;
  assign T_44456 = T_44455 & T_4324_94;
  assign T_44457 = T_44456 & T_4324_93;
  assign T_44458 = T_44457 & T_4324_92;
  assign T_44459 = T_44458 & T_4324_91;
  assign T_44460 = T_44459 & T_4324_90;
  assign T_44461 = T_44460 & T_4324_89;
  assign T_44462 = T_44461 & T_4324_88;
  assign T_44463 = T_44462 & T_4324_87;
  assign T_44464 = T_44463 & T_4324_86;
  assign T_44465 = T_44464 & T_4324_85;
  assign T_44466 = T_44465 & T_4324_84;
  assign T_44467 = T_44466 & T_4324_83;
  assign T_44468 = T_44467 & T_4324_82;
  assign T_44469 = T_44468 & T_4324_81;
  assign T_44470 = T_44469 & T_4324_80;
  assign T_44471 = T_44470 & T_4324_79;
  assign T_44480 = T_41407 & T_4329_102;
  assign T_44481 = T_44480 & T_4329_101;
  assign T_44482 = T_44481 & T_4329_100;
  assign T_44483 = T_44482 & T_4329_99;
  assign T_44484 = T_44483 & T_4329_98;
  assign T_44485 = T_44484 & T_4329_97;
  assign T_44486 = T_44485 & T_4329_96;
  assign T_44487 = T_44486 & T_4329_95;
  assign T_44488 = T_44487 & T_4329_94;
  assign T_44489 = T_44488 & T_4329_93;
  assign T_44490 = T_44489 & T_4329_92;
  assign T_44491 = T_44490 & T_4329_91;
  assign T_44492 = T_44491 & T_4329_90;
  assign T_44493 = T_44492 & T_4329_89;
  assign T_44494 = T_44493 & T_4329_88;
  assign T_44495 = T_44494 & T_4329_87;
  assign T_44496 = T_44495 & T_4329_86;
  assign T_44497 = T_44496 & T_4329_85;
  assign T_44498 = T_44497 & T_4329_84;
  assign T_44499 = T_44498 & T_4329_83;
  assign T_44500 = T_44499 & T_4329_82;
  assign T_44501 = T_44500 & T_4329_81;
  assign T_44502 = T_44501 & T_4329_80;
  assign T_44503 = T_44502 & T_4329_79;
  assign T_44512 = T_41439 & T_4334_102;
  assign T_44513 = T_44512 & T_4334_101;
  assign T_44514 = T_44513 & T_4334_100;
  assign T_44515 = T_44514 & T_4334_99;
  assign T_44516 = T_44515 & T_4334_98;
  assign T_44517 = T_44516 & T_4334_97;
  assign T_44518 = T_44517 & T_4334_96;
  assign T_44519 = T_44518 & T_4334_95;
  assign T_44520 = T_44519 & T_4334_94;
  assign T_44521 = T_44520 & T_4334_93;
  assign T_44522 = T_44521 & T_4334_92;
  assign T_44523 = T_44522 & T_4334_91;
  assign T_44524 = T_44523 & T_4334_90;
  assign T_44525 = T_44524 & T_4334_89;
  assign T_44526 = T_44525 & T_4334_88;
  assign T_44527 = T_44526 & T_4334_87;
  assign T_44528 = T_44527 & T_4334_86;
  assign T_44529 = T_44528 & T_4334_85;
  assign T_44530 = T_44529 & T_4334_84;
  assign T_44531 = T_44530 & T_4334_83;
  assign T_44532 = T_44531 & T_4334_82;
  assign T_44533 = T_44532 & T_4334_81;
  assign T_44534 = T_44533 & T_4334_80;
  assign T_44535 = T_44534 & T_4334_79;
  assign T_44543 = T_41342 & T_4319_103;
  assign T_44544 = T_44543 & T_4319_102;
  assign T_44545 = T_44544 & T_4319_101;
  assign T_44546 = T_44545 & T_4319_100;
  assign T_44547 = T_44546 & T_4319_99;
  assign T_44548 = T_44547 & T_4319_98;
  assign T_44549 = T_44548 & T_4319_97;
  assign T_44550 = T_44549 & T_4319_96;
  assign T_44551 = T_44550 & T_4319_95;
  assign T_44552 = T_44551 & T_4319_94;
  assign T_44553 = T_44552 & T_4319_93;
  assign T_44554 = T_44553 & T_4319_92;
  assign T_44555 = T_44554 & T_4319_91;
  assign T_44556 = T_44555 & T_4319_90;
  assign T_44557 = T_44556 & T_4319_89;
  assign T_44558 = T_44557 & T_4319_88;
  assign T_44559 = T_44558 & T_4319_87;
  assign T_44560 = T_44559 & T_4319_86;
  assign T_44561 = T_44560 & T_4319_85;
  assign T_44562 = T_44561 & T_4319_84;
  assign T_44563 = T_44562 & T_4319_83;
  assign T_44564 = T_44563 & T_4319_82;
  assign T_44565 = T_44564 & T_4319_81;
  assign T_44566 = T_44565 & T_4319_80;
  assign T_44567 = T_44566 & T_4319_79;
  assign T_44575 = T_41374 & T_4324_103;
  assign T_44576 = T_44575 & T_4324_102;
  assign T_44577 = T_44576 & T_4324_101;
  assign T_44578 = T_44577 & T_4324_100;
  assign T_44579 = T_44578 & T_4324_99;
  assign T_44580 = T_44579 & T_4324_98;
  assign T_44581 = T_44580 & T_4324_97;
  assign T_44582 = T_44581 & T_4324_96;
  assign T_44583 = T_44582 & T_4324_95;
  assign T_44584 = T_44583 & T_4324_94;
  assign T_44585 = T_44584 & T_4324_93;
  assign T_44586 = T_44585 & T_4324_92;
  assign T_44587 = T_44586 & T_4324_91;
  assign T_44588 = T_44587 & T_4324_90;
  assign T_44589 = T_44588 & T_4324_89;
  assign T_44590 = T_44589 & T_4324_88;
  assign T_44591 = T_44590 & T_4324_87;
  assign T_44592 = T_44591 & T_4324_86;
  assign T_44593 = T_44592 & T_4324_85;
  assign T_44594 = T_44593 & T_4324_84;
  assign T_44595 = T_44594 & T_4324_83;
  assign T_44596 = T_44595 & T_4324_82;
  assign T_44597 = T_44596 & T_4324_81;
  assign T_44598 = T_44597 & T_4324_80;
  assign T_44599 = T_44598 & T_4324_79;
  assign T_44607 = T_41406 & T_4329_103;
  assign T_44608 = T_44607 & T_4329_102;
  assign T_44609 = T_44608 & T_4329_101;
  assign T_44610 = T_44609 & T_4329_100;
  assign T_44611 = T_44610 & T_4329_99;
  assign T_44612 = T_44611 & T_4329_98;
  assign T_44613 = T_44612 & T_4329_97;
  assign T_44614 = T_44613 & T_4329_96;
  assign T_44615 = T_44614 & T_4329_95;
  assign T_44616 = T_44615 & T_4329_94;
  assign T_44617 = T_44616 & T_4329_93;
  assign T_44618 = T_44617 & T_4329_92;
  assign T_44619 = T_44618 & T_4329_91;
  assign T_44620 = T_44619 & T_4329_90;
  assign T_44621 = T_44620 & T_4329_89;
  assign T_44622 = T_44621 & T_4329_88;
  assign T_44623 = T_44622 & T_4329_87;
  assign T_44624 = T_44623 & T_4329_86;
  assign T_44625 = T_44624 & T_4329_85;
  assign T_44626 = T_44625 & T_4329_84;
  assign T_44627 = T_44626 & T_4329_83;
  assign T_44628 = T_44627 & T_4329_82;
  assign T_44629 = T_44628 & T_4329_81;
  assign T_44630 = T_44629 & T_4329_80;
  assign T_44631 = T_44630 & T_4329_79;
  assign T_44639 = T_41438 & T_4334_103;
  assign T_44640 = T_44639 & T_4334_102;
  assign T_44641 = T_44640 & T_4334_101;
  assign T_44642 = T_44641 & T_4334_100;
  assign T_44643 = T_44642 & T_4334_99;
  assign T_44644 = T_44643 & T_4334_98;
  assign T_44645 = T_44644 & T_4334_97;
  assign T_44646 = T_44645 & T_4334_96;
  assign T_44647 = T_44646 & T_4334_95;
  assign T_44648 = T_44647 & T_4334_94;
  assign T_44649 = T_44648 & T_4334_93;
  assign T_44650 = T_44649 & T_4334_92;
  assign T_44651 = T_44650 & T_4334_91;
  assign T_44652 = T_44651 & T_4334_90;
  assign T_44653 = T_44652 & T_4334_89;
  assign T_44654 = T_44653 & T_4334_88;
  assign T_44655 = T_44654 & T_4334_87;
  assign T_44656 = T_44655 & T_4334_86;
  assign T_44657 = T_44656 & T_4334_85;
  assign T_44658 = T_44657 & T_4334_84;
  assign T_44659 = T_44658 & T_4334_83;
  assign T_44660 = T_44659 & T_4334_82;
  assign T_44661 = T_44660 & T_4334_81;
  assign T_44662 = T_44661 & T_4334_80;
  assign T_44663 = T_44662 & T_4334_79;
  assign T_44670 = T_41341 & T_4319_104;
  assign T_44671 = T_44670 & T_4319_103;
  assign T_44672 = T_44671 & T_4319_102;
  assign T_44673 = T_44672 & T_4319_101;
  assign T_44674 = T_44673 & T_4319_100;
  assign T_44675 = T_44674 & T_4319_99;
  assign T_44676 = T_44675 & T_4319_98;
  assign T_44677 = T_44676 & T_4319_97;
  assign T_44678 = T_44677 & T_4319_96;
  assign T_44679 = T_44678 & T_4319_95;
  assign T_44680 = T_44679 & T_4319_94;
  assign T_44681 = T_44680 & T_4319_93;
  assign T_44682 = T_44681 & T_4319_92;
  assign T_44683 = T_44682 & T_4319_91;
  assign T_44684 = T_44683 & T_4319_90;
  assign T_44685 = T_44684 & T_4319_89;
  assign T_44686 = T_44685 & T_4319_88;
  assign T_44687 = T_44686 & T_4319_87;
  assign T_44688 = T_44687 & T_4319_86;
  assign T_44689 = T_44688 & T_4319_85;
  assign T_44690 = T_44689 & T_4319_84;
  assign T_44691 = T_44690 & T_4319_83;
  assign T_44692 = T_44691 & T_4319_82;
  assign T_44693 = T_44692 & T_4319_81;
  assign T_44694 = T_44693 & T_4319_80;
  assign T_44695 = T_44694 & T_4319_79;
  assign T_44702 = T_41373 & T_4324_104;
  assign T_44703 = T_44702 & T_4324_103;
  assign T_44704 = T_44703 & T_4324_102;
  assign T_44705 = T_44704 & T_4324_101;
  assign T_44706 = T_44705 & T_4324_100;
  assign T_44707 = T_44706 & T_4324_99;
  assign T_44708 = T_44707 & T_4324_98;
  assign T_44709 = T_44708 & T_4324_97;
  assign T_44710 = T_44709 & T_4324_96;
  assign T_44711 = T_44710 & T_4324_95;
  assign T_44712 = T_44711 & T_4324_94;
  assign T_44713 = T_44712 & T_4324_93;
  assign T_44714 = T_44713 & T_4324_92;
  assign T_44715 = T_44714 & T_4324_91;
  assign T_44716 = T_44715 & T_4324_90;
  assign T_44717 = T_44716 & T_4324_89;
  assign T_44718 = T_44717 & T_4324_88;
  assign T_44719 = T_44718 & T_4324_87;
  assign T_44720 = T_44719 & T_4324_86;
  assign T_44721 = T_44720 & T_4324_85;
  assign T_44722 = T_44721 & T_4324_84;
  assign T_44723 = T_44722 & T_4324_83;
  assign T_44724 = T_44723 & T_4324_82;
  assign T_44725 = T_44724 & T_4324_81;
  assign T_44726 = T_44725 & T_4324_80;
  assign T_44727 = T_44726 & T_4324_79;
  assign T_44734 = T_41405 & T_4329_104;
  assign T_44735 = T_44734 & T_4329_103;
  assign T_44736 = T_44735 & T_4329_102;
  assign T_44737 = T_44736 & T_4329_101;
  assign T_44738 = T_44737 & T_4329_100;
  assign T_44739 = T_44738 & T_4329_99;
  assign T_44740 = T_44739 & T_4329_98;
  assign T_44741 = T_44740 & T_4329_97;
  assign T_44742 = T_44741 & T_4329_96;
  assign T_44743 = T_44742 & T_4329_95;
  assign T_44744 = T_44743 & T_4329_94;
  assign T_44745 = T_44744 & T_4329_93;
  assign T_44746 = T_44745 & T_4329_92;
  assign T_44747 = T_44746 & T_4329_91;
  assign T_44748 = T_44747 & T_4329_90;
  assign T_44749 = T_44748 & T_4329_89;
  assign T_44750 = T_44749 & T_4329_88;
  assign T_44751 = T_44750 & T_4329_87;
  assign T_44752 = T_44751 & T_4329_86;
  assign T_44753 = T_44752 & T_4329_85;
  assign T_44754 = T_44753 & T_4329_84;
  assign T_44755 = T_44754 & T_4329_83;
  assign T_44756 = T_44755 & T_4329_82;
  assign T_44757 = T_44756 & T_4329_81;
  assign T_44758 = T_44757 & T_4329_80;
  assign T_44759 = T_44758 & T_4329_79;
  assign T_44766 = T_41437 & T_4334_104;
  assign T_44767 = T_44766 & T_4334_103;
  assign T_44768 = T_44767 & T_4334_102;
  assign T_44769 = T_44768 & T_4334_101;
  assign T_44770 = T_44769 & T_4334_100;
  assign T_44771 = T_44770 & T_4334_99;
  assign T_44772 = T_44771 & T_4334_98;
  assign T_44773 = T_44772 & T_4334_97;
  assign T_44774 = T_44773 & T_4334_96;
  assign T_44775 = T_44774 & T_4334_95;
  assign T_44776 = T_44775 & T_4334_94;
  assign T_44777 = T_44776 & T_4334_93;
  assign T_44778 = T_44777 & T_4334_92;
  assign T_44779 = T_44778 & T_4334_91;
  assign T_44780 = T_44779 & T_4334_90;
  assign T_44781 = T_44780 & T_4334_89;
  assign T_44782 = T_44781 & T_4334_88;
  assign T_44783 = T_44782 & T_4334_87;
  assign T_44784 = T_44783 & T_4334_86;
  assign T_44785 = T_44784 & T_4334_85;
  assign T_44786 = T_44785 & T_4334_84;
  assign T_44787 = T_44786 & T_4334_83;
  assign T_44788 = T_44787 & T_4334_82;
  assign T_44789 = T_44788 & T_4334_81;
  assign T_44790 = T_44789 & T_4334_80;
  assign T_44791 = T_44790 & T_4334_79;
  assign T_44797 = T_41340 & T_4319_105;
  assign T_44798 = T_44797 & T_4319_104;
  assign T_44799 = T_44798 & T_4319_103;
  assign T_44800 = T_44799 & T_4319_102;
  assign T_44801 = T_44800 & T_4319_101;
  assign T_44802 = T_44801 & T_4319_100;
  assign T_44803 = T_44802 & T_4319_99;
  assign T_44804 = T_44803 & T_4319_98;
  assign T_44805 = T_44804 & T_4319_97;
  assign T_44806 = T_44805 & T_4319_96;
  assign T_44807 = T_44806 & T_4319_95;
  assign T_44808 = T_44807 & T_4319_94;
  assign T_44809 = T_44808 & T_4319_93;
  assign T_44810 = T_44809 & T_4319_92;
  assign T_44811 = T_44810 & T_4319_91;
  assign T_44812 = T_44811 & T_4319_90;
  assign T_44813 = T_44812 & T_4319_89;
  assign T_44814 = T_44813 & T_4319_88;
  assign T_44815 = T_44814 & T_4319_87;
  assign T_44816 = T_44815 & T_4319_86;
  assign T_44817 = T_44816 & T_4319_85;
  assign T_44818 = T_44817 & T_4319_84;
  assign T_44819 = T_44818 & T_4319_83;
  assign T_44820 = T_44819 & T_4319_82;
  assign T_44821 = T_44820 & T_4319_81;
  assign T_44822 = T_44821 & T_4319_80;
  assign T_44823 = T_44822 & T_4319_79;
  assign T_44829 = T_41372 & T_4324_105;
  assign T_44830 = T_44829 & T_4324_104;
  assign T_44831 = T_44830 & T_4324_103;
  assign T_44832 = T_44831 & T_4324_102;
  assign T_44833 = T_44832 & T_4324_101;
  assign T_44834 = T_44833 & T_4324_100;
  assign T_44835 = T_44834 & T_4324_99;
  assign T_44836 = T_44835 & T_4324_98;
  assign T_44837 = T_44836 & T_4324_97;
  assign T_44838 = T_44837 & T_4324_96;
  assign T_44839 = T_44838 & T_4324_95;
  assign T_44840 = T_44839 & T_4324_94;
  assign T_44841 = T_44840 & T_4324_93;
  assign T_44842 = T_44841 & T_4324_92;
  assign T_44843 = T_44842 & T_4324_91;
  assign T_44844 = T_44843 & T_4324_90;
  assign T_44845 = T_44844 & T_4324_89;
  assign T_44846 = T_44845 & T_4324_88;
  assign T_44847 = T_44846 & T_4324_87;
  assign T_44848 = T_44847 & T_4324_86;
  assign T_44849 = T_44848 & T_4324_85;
  assign T_44850 = T_44849 & T_4324_84;
  assign T_44851 = T_44850 & T_4324_83;
  assign T_44852 = T_44851 & T_4324_82;
  assign T_44853 = T_44852 & T_4324_81;
  assign T_44854 = T_44853 & T_4324_80;
  assign T_44855 = T_44854 & T_4324_79;
  assign T_44861 = T_41404 & T_4329_105;
  assign T_44862 = T_44861 & T_4329_104;
  assign T_44863 = T_44862 & T_4329_103;
  assign T_44864 = T_44863 & T_4329_102;
  assign T_44865 = T_44864 & T_4329_101;
  assign T_44866 = T_44865 & T_4329_100;
  assign T_44867 = T_44866 & T_4329_99;
  assign T_44868 = T_44867 & T_4329_98;
  assign T_44869 = T_44868 & T_4329_97;
  assign T_44870 = T_44869 & T_4329_96;
  assign T_44871 = T_44870 & T_4329_95;
  assign T_44872 = T_44871 & T_4329_94;
  assign T_44873 = T_44872 & T_4329_93;
  assign T_44874 = T_44873 & T_4329_92;
  assign T_44875 = T_44874 & T_4329_91;
  assign T_44876 = T_44875 & T_4329_90;
  assign T_44877 = T_44876 & T_4329_89;
  assign T_44878 = T_44877 & T_4329_88;
  assign T_44879 = T_44878 & T_4329_87;
  assign T_44880 = T_44879 & T_4329_86;
  assign T_44881 = T_44880 & T_4329_85;
  assign T_44882 = T_44881 & T_4329_84;
  assign T_44883 = T_44882 & T_4329_83;
  assign T_44884 = T_44883 & T_4329_82;
  assign T_44885 = T_44884 & T_4329_81;
  assign T_44886 = T_44885 & T_4329_80;
  assign T_44887 = T_44886 & T_4329_79;
  assign T_44893 = T_41436 & T_4334_105;
  assign T_44894 = T_44893 & T_4334_104;
  assign T_44895 = T_44894 & T_4334_103;
  assign T_44896 = T_44895 & T_4334_102;
  assign T_44897 = T_44896 & T_4334_101;
  assign T_44898 = T_44897 & T_4334_100;
  assign T_44899 = T_44898 & T_4334_99;
  assign T_44900 = T_44899 & T_4334_98;
  assign T_44901 = T_44900 & T_4334_97;
  assign T_44902 = T_44901 & T_4334_96;
  assign T_44903 = T_44902 & T_4334_95;
  assign T_44904 = T_44903 & T_4334_94;
  assign T_44905 = T_44904 & T_4334_93;
  assign T_44906 = T_44905 & T_4334_92;
  assign T_44907 = T_44906 & T_4334_91;
  assign T_44908 = T_44907 & T_4334_90;
  assign T_44909 = T_44908 & T_4334_89;
  assign T_44910 = T_44909 & T_4334_88;
  assign T_44911 = T_44910 & T_4334_87;
  assign T_44912 = T_44911 & T_4334_86;
  assign T_44913 = T_44912 & T_4334_85;
  assign T_44914 = T_44913 & T_4334_84;
  assign T_44915 = T_44914 & T_4334_83;
  assign T_44916 = T_44915 & T_4334_82;
  assign T_44917 = T_44916 & T_4334_81;
  assign T_44918 = T_44917 & T_4334_80;
  assign T_44919 = T_44918 & T_4334_79;
  assign T_44924 = T_41339 & T_4319_106;
  assign T_44925 = T_44924 & T_4319_105;
  assign T_44926 = T_44925 & T_4319_104;
  assign T_44927 = T_44926 & T_4319_103;
  assign T_44928 = T_44927 & T_4319_102;
  assign T_44929 = T_44928 & T_4319_101;
  assign T_44930 = T_44929 & T_4319_100;
  assign T_44931 = T_44930 & T_4319_99;
  assign T_44932 = T_44931 & T_4319_98;
  assign T_44933 = T_44932 & T_4319_97;
  assign T_44934 = T_44933 & T_4319_96;
  assign T_44935 = T_44934 & T_4319_95;
  assign T_44936 = T_44935 & T_4319_94;
  assign T_44937 = T_44936 & T_4319_93;
  assign T_44938 = T_44937 & T_4319_92;
  assign T_44939 = T_44938 & T_4319_91;
  assign T_44940 = T_44939 & T_4319_90;
  assign T_44941 = T_44940 & T_4319_89;
  assign T_44942 = T_44941 & T_4319_88;
  assign T_44943 = T_44942 & T_4319_87;
  assign T_44944 = T_44943 & T_4319_86;
  assign T_44945 = T_44944 & T_4319_85;
  assign T_44946 = T_44945 & T_4319_84;
  assign T_44947 = T_44946 & T_4319_83;
  assign T_44948 = T_44947 & T_4319_82;
  assign T_44949 = T_44948 & T_4319_81;
  assign T_44950 = T_44949 & T_4319_80;
  assign T_44951 = T_44950 & T_4319_79;
  assign T_44956 = T_41371 & T_4324_106;
  assign T_44957 = T_44956 & T_4324_105;
  assign T_44958 = T_44957 & T_4324_104;
  assign T_44959 = T_44958 & T_4324_103;
  assign T_44960 = T_44959 & T_4324_102;
  assign T_44961 = T_44960 & T_4324_101;
  assign T_44962 = T_44961 & T_4324_100;
  assign T_44963 = T_44962 & T_4324_99;
  assign T_44964 = T_44963 & T_4324_98;
  assign T_44965 = T_44964 & T_4324_97;
  assign T_44966 = T_44965 & T_4324_96;
  assign T_44967 = T_44966 & T_4324_95;
  assign T_44968 = T_44967 & T_4324_94;
  assign T_44969 = T_44968 & T_4324_93;
  assign T_44970 = T_44969 & T_4324_92;
  assign T_44971 = T_44970 & T_4324_91;
  assign T_44972 = T_44971 & T_4324_90;
  assign T_44973 = T_44972 & T_4324_89;
  assign T_44974 = T_44973 & T_4324_88;
  assign T_44975 = T_44974 & T_4324_87;
  assign T_44976 = T_44975 & T_4324_86;
  assign T_44977 = T_44976 & T_4324_85;
  assign T_44978 = T_44977 & T_4324_84;
  assign T_44979 = T_44978 & T_4324_83;
  assign T_44980 = T_44979 & T_4324_82;
  assign T_44981 = T_44980 & T_4324_81;
  assign T_44982 = T_44981 & T_4324_80;
  assign T_44983 = T_44982 & T_4324_79;
  assign T_44988 = T_41403 & T_4329_106;
  assign T_44989 = T_44988 & T_4329_105;
  assign T_44990 = T_44989 & T_4329_104;
  assign T_44991 = T_44990 & T_4329_103;
  assign T_44992 = T_44991 & T_4329_102;
  assign T_44993 = T_44992 & T_4329_101;
  assign T_44994 = T_44993 & T_4329_100;
  assign T_44995 = T_44994 & T_4329_99;
  assign T_44996 = T_44995 & T_4329_98;
  assign T_44997 = T_44996 & T_4329_97;
  assign T_44998 = T_44997 & T_4329_96;
  assign T_44999 = T_44998 & T_4329_95;
  assign T_45000 = T_44999 & T_4329_94;
  assign T_45001 = T_45000 & T_4329_93;
  assign T_45002 = T_45001 & T_4329_92;
  assign T_45003 = T_45002 & T_4329_91;
  assign T_45004 = T_45003 & T_4329_90;
  assign T_45005 = T_45004 & T_4329_89;
  assign T_45006 = T_45005 & T_4329_88;
  assign T_45007 = T_45006 & T_4329_87;
  assign T_45008 = T_45007 & T_4329_86;
  assign T_45009 = T_45008 & T_4329_85;
  assign T_45010 = T_45009 & T_4329_84;
  assign T_45011 = T_45010 & T_4329_83;
  assign T_45012 = T_45011 & T_4329_82;
  assign T_45013 = T_45012 & T_4329_81;
  assign T_45014 = T_45013 & T_4329_80;
  assign T_45015 = T_45014 & T_4329_79;
  assign T_45020 = T_41435 & T_4334_106;
  assign T_45021 = T_45020 & T_4334_105;
  assign T_45022 = T_45021 & T_4334_104;
  assign T_45023 = T_45022 & T_4334_103;
  assign T_45024 = T_45023 & T_4334_102;
  assign T_45025 = T_45024 & T_4334_101;
  assign T_45026 = T_45025 & T_4334_100;
  assign T_45027 = T_45026 & T_4334_99;
  assign T_45028 = T_45027 & T_4334_98;
  assign T_45029 = T_45028 & T_4334_97;
  assign T_45030 = T_45029 & T_4334_96;
  assign T_45031 = T_45030 & T_4334_95;
  assign T_45032 = T_45031 & T_4334_94;
  assign T_45033 = T_45032 & T_4334_93;
  assign T_45034 = T_45033 & T_4334_92;
  assign T_45035 = T_45034 & T_4334_91;
  assign T_45036 = T_45035 & T_4334_90;
  assign T_45037 = T_45036 & T_4334_89;
  assign T_45038 = T_45037 & T_4334_88;
  assign T_45039 = T_45038 & T_4334_87;
  assign T_45040 = T_45039 & T_4334_86;
  assign T_45041 = T_45040 & T_4334_85;
  assign T_45042 = T_45041 & T_4334_84;
  assign T_45043 = T_45042 & T_4334_83;
  assign T_45044 = T_45043 & T_4334_82;
  assign T_45045 = T_45044 & T_4334_81;
  assign T_45046 = T_45045 & T_4334_80;
  assign T_45047 = T_45046 & T_4334_79;
  assign T_45051 = T_41338 & T_4319_107;
  assign T_45052 = T_45051 & T_4319_106;
  assign T_45053 = T_45052 & T_4319_105;
  assign T_45054 = T_45053 & T_4319_104;
  assign T_45055 = T_45054 & T_4319_103;
  assign T_45056 = T_45055 & T_4319_102;
  assign T_45057 = T_45056 & T_4319_101;
  assign T_45058 = T_45057 & T_4319_100;
  assign T_45059 = T_45058 & T_4319_99;
  assign T_45060 = T_45059 & T_4319_98;
  assign T_45061 = T_45060 & T_4319_97;
  assign T_45062 = T_45061 & T_4319_96;
  assign T_45063 = T_45062 & T_4319_95;
  assign T_45064 = T_45063 & T_4319_94;
  assign T_45065 = T_45064 & T_4319_93;
  assign T_45066 = T_45065 & T_4319_92;
  assign T_45067 = T_45066 & T_4319_91;
  assign T_45068 = T_45067 & T_4319_90;
  assign T_45069 = T_45068 & T_4319_89;
  assign T_45070 = T_45069 & T_4319_88;
  assign T_45071 = T_45070 & T_4319_87;
  assign T_45072 = T_45071 & T_4319_86;
  assign T_45073 = T_45072 & T_4319_85;
  assign T_45074 = T_45073 & T_4319_84;
  assign T_45075 = T_45074 & T_4319_83;
  assign T_45076 = T_45075 & T_4319_82;
  assign T_45077 = T_45076 & T_4319_81;
  assign T_45078 = T_45077 & T_4319_80;
  assign T_45079 = T_45078 & T_4319_79;
  assign T_45083 = T_41370 & T_4324_107;
  assign T_45084 = T_45083 & T_4324_106;
  assign T_45085 = T_45084 & T_4324_105;
  assign T_45086 = T_45085 & T_4324_104;
  assign T_45087 = T_45086 & T_4324_103;
  assign T_45088 = T_45087 & T_4324_102;
  assign T_45089 = T_45088 & T_4324_101;
  assign T_45090 = T_45089 & T_4324_100;
  assign T_45091 = T_45090 & T_4324_99;
  assign T_45092 = T_45091 & T_4324_98;
  assign T_45093 = T_45092 & T_4324_97;
  assign T_45094 = T_45093 & T_4324_96;
  assign T_45095 = T_45094 & T_4324_95;
  assign T_45096 = T_45095 & T_4324_94;
  assign T_45097 = T_45096 & T_4324_93;
  assign T_45098 = T_45097 & T_4324_92;
  assign T_45099 = T_45098 & T_4324_91;
  assign T_45100 = T_45099 & T_4324_90;
  assign T_45101 = T_45100 & T_4324_89;
  assign T_45102 = T_45101 & T_4324_88;
  assign T_45103 = T_45102 & T_4324_87;
  assign T_45104 = T_45103 & T_4324_86;
  assign T_45105 = T_45104 & T_4324_85;
  assign T_45106 = T_45105 & T_4324_84;
  assign T_45107 = T_45106 & T_4324_83;
  assign T_45108 = T_45107 & T_4324_82;
  assign T_45109 = T_45108 & T_4324_81;
  assign T_45110 = T_45109 & T_4324_80;
  assign T_45111 = T_45110 & T_4324_79;
  assign T_45115 = T_41402 & T_4329_107;
  assign T_45116 = T_45115 & T_4329_106;
  assign T_45117 = T_45116 & T_4329_105;
  assign T_45118 = T_45117 & T_4329_104;
  assign T_45119 = T_45118 & T_4329_103;
  assign T_45120 = T_45119 & T_4329_102;
  assign T_45121 = T_45120 & T_4329_101;
  assign T_45122 = T_45121 & T_4329_100;
  assign T_45123 = T_45122 & T_4329_99;
  assign T_45124 = T_45123 & T_4329_98;
  assign T_45125 = T_45124 & T_4329_97;
  assign T_45126 = T_45125 & T_4329_96;
  assign T_45127 = T_45126 & T_4329_95;
  assign T_45128 = T_45127 & T_4329_94;
  assign T_45129 = T_45128 & T_4329_93;
  assign T_45130 = T_45129 & T_4329_92;
  assign T_45131 = T_45130 & T_4329_91;
  assign T_45132 = T_45131 & T_4329_90;
  assign T_45133 = T_45132 & T_4329_89;
  assign T_45134 = T_45133 & T_4329_88;
  assign T_45135 = T_45134 & T_4329_87;
  assign T_45136 = T_45135 & T_4329_86;
  assign T_45137 = T_45136 & T_4329_85;
  assign T_45138 = T_45137 & T_4329_84;
  assign T_45139 = T_45138 & T_4329_83;
  assign T_45140 = T_45139 & T_4329_82;
  assign T_45141 = T_45140 & T_4329_81;
  assign T_45142 = T_45141 & T_4329_80;
  assign T_45143 = T_45142 & T_4329_79;
  assign T_45147 = T_41434 & T_4334_107;
  assign T_45148 = T_45147 & T_4334_106;
  assign T_45149 = T_45148 & T_4334_105;
  assign T_45150 = T_45149 & T_4334_104;
  assign T_45151 = T_45150 & T_4334_103;
  assign T_45152 = T_45151 & T_4334_102;
  assign T_45153 = T_45152 & T_4334_101;
  assign T_45154 = T_45153 & T_4334_100;
  assign T_45155 = T_45154 & T_4334_99;
  assign T_45156 = T_45155 & T_4334_98;
  assign T_45157 = T_45156 & T_4334_97;
  assign T_45158 = T_45157 & T_4334_96;
  assign T_45159 = T_45158 & T_4334_95;
  assign T_45160 = T_45159 & T_4334_94;
  assign T_45161 = T_45160 & T_4334_93;
  assign T_45162 = T_45161 & T_4334_92;
  assign T_45163 = T_45162 & T_4334_91;
  assign T_45164 = T_45163 & T_4334_90;
  assign T_45165 = T_45164 & T_4334_89;
  assign T_45166 = T_45165 & T_4334_88;
  assign T_45167 = T_45166 & T_4334_87;
  assign T_45168 = T_45167 & T_4334_86;
  assign T_45169 = T_45168 & T_4334_85;
  assign T_45170 = T_45169 & T_4334_84;
  assign T_45171 = T_45170 & T_4334_83;
  assign T_45172 = T_45171 & T_4334_82;
  assign T_45173 = T_45172 & T_4334_81;
  assign T_45174 = T_45173 & T_4334_80;
  assign T_45175 = T_45174 & T_4334_79;
  assign T_45178 = T_41337 & T_4319_108;
  assign T_45179 = T_45178 & T_4319_107;
  assign T_45180 = T_45179 & T_4319_106;
  assign T_45181 = T_45180 & T_4319_105;
  assign T_45182 = T_45181 & T_4319_104;
  assign T_45183 = T_45182 & T_4319_103;
  assign T_45184 = T_45183 & T_4319_102;
  assign T_45185 = T_45184 & T_4319_101;
  assign T_45186 = T_45185 & T_4319_100;
  assign T_45187 = T_45186 & T_4319_99;
  assign T_45188 = T_45187 & T_4319_98;
  assign T_45189 = T_45188 & T_4319_97;
  assign T_45190 = T_45189 & T_4319_96;
  assign T_45191 = T_45190 & T_4319_95;
  assign T_45192 = T_45191 & T_4319_94;
  assign T_45193 = T_45192 & T_4319_93;
  assign T_45194 = T_45193 & T_4319_92;
  assign T_45195 = T_45194 & T_4319_91;
  assign T_45196 = T_45195 & T_4319_90;
  assign T_45197 = T_45196 & T_4319_89;
  assign T_45198 = T_45197 & T_4319_88;
  assign T_45199 = T_45198 & T_4319_87;
  assign T_45200 = T_45199 & T_4319_86;
  assign T_45201 = T_45200 & T_4319_85;
  assign T_45202 = T_45201 & T_4319_84;
  assign T_45203 = T_45202 & T_4319_83;
  assign T_45204 = T_45203 & T_4319_82;
  assign T_45205 = T_45204 & T_4319_81;
  assign T_45206 = T_45205 & T_4319_80;
  assign T_45207 = T_45206 & T_4319_79;
  assign T_45210 = T_41369 & T_4324_108;
  assign T_45211 = T_45210 & T_4324_107;
  assign T_45212 = T_45211 & T_4324_106;
  assign T_45213 = T_45212 & T_4324_105;
  assign T_45214 = T_45213 & T_4324_104;
  assign T_45215 = T_45214 & T_4324_103;
  assign T_45216 = T_45215 & T_4324_102;
  assign T_45217 = T_45216 & T_4324_101;
  assign T_45218 = T_45217 & T_4324_100;
  assign T_45219 = T_45218 & T_4324_99;
  assign T_45220 = T_45219 & T_4324_98;
  assign T_45221 = T_45220 & T_4324_97;
  assign T_45222 = T_45221 & T_4324_96;
  assign T_45223 = T_45222 & T_4324_95;
  assign T_45224 = T_45223 & T_4324_94;
  assign T_45225 = T_45224 & T_4324_93;
  assign T_45226 = T_45225 & T_4324_92;
  assign T_45227 = T_45226 & T_4324_91;
  assign T_45228 = T_45227 & T_4324_90;
  assign T_45229 = T_45228 & T_4324_89;
  assign T_45230 = T_45229 & T_4324_88;
  assign T_45231 = T_45230 & T_4324_87;
  assign T_45232 = T_45231 & T_4324_86;
  assign T_45233 = T_45232 & T_4324_85;
  assign T_45234 = T_45233 & T_4324_84;
  assign T_45235 = T_45234 & T_4324_83;
  assign T_45236 = T_45235 & T_4324_82;
  assign T_45237 = T_45236 & T_4324_81;
  assign T_45238 = T_45237 & T_4324_80;
  assign T_45239 = T_45238 & T_4324_79;
  assign T_45242 = T_41401 & T_4329_108;
  assign T_45243 = T_45242 & T_4329_107;
  assign T_45244 = T_45243 & T_4329_106;
  assign T_45245 = T_45244 & T_4329_105;
  assign T_45246 = T_45245 & T_4329_104;
  assign T_45247 = T_45246 & T_4329_103;
  assign T_45248 = T_45247 & T_4329_102;
  assign T_45249 = T_45248 & T_4329_101;
  assign T_45250 = T_45249 & T_4329_100;
  assign T_45251 = T_45250 & T_4329_99;
  assign T_45252 = T_45251 & T_4329_98;
  assign T_45253 = T_45252 & T_4329_97;
  assign T_45254 = T_45253 & T_4329_96;
  assign T_45255 = T_45254 & T_4329_95;
  assign T_45256 = T_45255 & T_4329_94;
  assign T_45257 = T_45256 & T_4329_93;
  assign T_45258 = T_45257 & T_4329_92;
  assign T_45259 = T_45258 & T_4329_91;
  assign T_45260 = T_45259 & T_4329_90;
  assign T_45261 = T_45260 & T_4329_89;
  assign T_45262 = T_45261 & T_4329_88;
  assign T_45263 = T_45262 & T_4329_87;
  assign T_45264 = T_45263 & T_4329_86;
  assign T_45265 = T_45264 & T_4329_85;
  assign T_45266 = T_45265 & T_4329_84;
  assign T_45267 = T_45266 & T_4329_83;
  assign T_45268 = T_45267 & T_4329_82;
  assign T_45269 = T_45268 & T_4329_81;
  assign T_45270 = T_45269 & T_4329_80;
  assign T_45271 = T_45270 & T_4329_79;
  assign T_45274 = T_41433 & T_4334_108;
  assign T_45275 = T_45274 & T_4334_107;
  assign T_45276 = T_45275 & T_4334_106;
  assign T_45277 = T_45276 & T_4334_105;
  assign T_45278 = T_45277 & T_4334_104;
  assign T_45279 = T_45278 & T_4334_103;
  assign T_45280 = T_45279 & T_4334_102;
  assign T_45281 = T_45280 & T_4334_101;
  assign T_45282 = T_45281 & T_4334_100;
  assign T_45283 = T_45282 & T_4334_99;
  assign T_45284 = T_45283 & T_4334_98;
  assign T_45285 = T_45284 & T_4334_97;
  assign T_45286 = T_45285 & T_4334_96;
  assign T_45287 = T_45286 & T_4334_95;
  assign T_45288 = T_45287 & T_4334_94;
  assign T_45289 = T_45288 & T_4334_93;
  assign T_45290 = T_45289 & T_4334_92;
  assign T_45291 = T_45290 & T_4334_91;
  assign T_45292 = T_45291 & T_4334_90;
  assign T_45293 = T_45292 & T_4334_89;
  assign T_45294 = T_45293 & T_4334_88;
  assign T_45295 = T_45294 & T_4334_87;
  assign T_45296 = T_45295 & T_4334_86;
  assign T_45297 = T_45296 & T_4334_85;
  assign T_45298 = T_45297 & T_4334_84;
  assign T_45299 = T_45298 & T_4334_83;
  assign T_45300 = T_45299 & T_4334_82;
  assign T_45301 = T_45300 & T_4334_81;
  assign T_45302 = T_45301 & T_4334_80;
  assign T_45303 = T_45302 & T_4334_79;
  assign T_45305 = T_27856 & T_4319_109;
  assign T_45306 = T_45305 & T_4319_108;
  assign T_45307 = T_45306 & T_4319_107;
  assign T_45308 = T_45307 & T_4319_106;
  assign T_45309 = T_45308 & T_4319_105;
  assign T_45310 = T_45309 & T_4319_104;
  assign T_45311 = T_45310 & T_4319_103;
  assign T_45312 = T_45311 & T_4319_102;
  assign T_45313 = T_45312 & T_4319_101;
  assign T_45314 = T_45313 & T_4319_100;
  assign T_45315 = T_45314 & T_4319_99;
  assign T_45316 = T_45315 & T_4319_98;
  assign T_45317 = T_45316 & T_4319_97;
  assign T_45318 = T_45317 & T_4319_96;
  assign T_45319 = T_45318 & T_4319_95;
  assign T_45320 = T_45319 & T_4319_94;
  assign T_45321 = T_45320 & T_4319_93;
  assign T_45322 = T_45321 & T_4319_92;
  assign T_45323 = T_45322 & T_4319_91;
  assign T_45324 = T_45323 & T_4319_90;
  assign T_45325 = T_45324 & T_4319_89;
  assign T_45326 = T_45325 & T_4319_88;
  assign T_45327 = T_45326 & T_4319_87;
  assign T_45328 = T_45327 & T_4319_86;
  assign T_45329 = T_45328 & T_4319_85;
  assign T_45330 = T_45329 & T_4319_84;
  assign T_45331 = T_45330 & T_4319_83;
  assign T_45332 = T_45331 & T_4319_82;
  assign T_45333 = T_45332 & T_4319_81;
  assign T_45334 = T_45333 & T_4319_80;
  assign T_45335 = T_45334 & T_4319_79;
  assign T_45337 = T_27862 & T_4324_109;
  assign T_45338 = T_45337 & T_4324_108;
  assign T_45339 = T_45338 & T_4324_107;
  assign T_45340 = T_45339 & T_4324_106;
  assign T_45341 = T_45340 & T_4324_105;
  assign T_45342 = T_45341 & T_4324_104;
  assign T_45343 = T_45342 & T_4324_103;
  assign T_45344 = T_45343 & T_4324_102;
  assign T_45345 = T_45344 & T_4324_101;
  assign T_45346 = T_45345 & T_4324_100;
  assign T_45347 = T_45346 & T_4324_99;
  assign T_45348 = T_45347 & T_4324_98;
  assign T_45349 = T_45348 & T_4324_97;
  assign T_45350 = T_45349 & T_4324_96;
  assign T_45351 = T_45350 & T_4324_95;
  assign T_45352 = T_45351 & T_4324_94;
  assign T_45353 = T_45352 & T_4324_93;
  assign T_45354 = T_45353 & T_4324_92;
  assign T_45355 = T_45354 & T_4324_91;
  assign T_45356 = T_45355 & T_4324_90;
  assign T_45357 = T_45356 & T_4324_89;
  assign T_45358 = T_45357 & T_4324_88;
  assign T_45359 = T_45358 & T_4324_87;
  assign T_45360 = T_45359 & T_4324_86;
  assign T_45361 = T_45360 & T_4324_85;
  assign T_45362 = T_45361 & T_4324_84;
  assign T_45363 = T_45362 & T_4324_83;
  assign T_45364 = T_45363 & T_4324_82;
  assign T_45365 = T_45364 & T_4324_81;
  assign T_45366 = T_45365 & T_4324_80;
  assign T_45367 = T_45366 & T_4324_79;
  assign T_45369 = T_27866 & T_4329_109;
  assign T_45370 = T_45369 & T_4329_108;
  assign T_45371 = T_45370 & T_4329_107;
  assign T_45372 = T_45371 & T_4329_106;
  assign T_45373 = T_45372 & T_4329_105;
  assign T_45374 = T_45373 & T_4329_104;
  assign T_45375 = T_45374 & T_4329_103;
  assign T_45376 = T_45375 & T_4329_102;
  assign T_45377 = T_45376 & T_4329_101;
  assign T_45378 = T_45377 & T_4329_100;
  assign T_45379 = T_45378 & T_4329_99;
  assign T_45380 = T_45379 & T_4329_98;
  assign T_45381 = T_45380 & T_4329_97;
  assign T_45382 = T_45381 & T_4329_96;
  assign T_45383 = T_45382 & T_4329_95;
  assign T_45384 = T_45383 & T_4329_94;
  assign T_45385 = T_45384 & T_4329_93;
  assign T_45386 = T_45385 & T_4329_92;
  assign T_45387 = T_45386 & T_4329_91;
  assign T_45388 = T_45387 & T_4329_90;
  assign T_45389 = T_45388 & T_4329_89;
  assign T_45390 = T_45389 & T_4329_88;
  assign T_45391 = T_45390 & T_4329_87;
  assign T_45392 = T_45391 & T_4329_86;
  assign T_45393 = T_45392 & T_4329_85;
  assign T_45394 = T_45393 & T_4329_84;
  assign T_45395 = T_45394 & T_4329_83;
  assign T_45396 = T_45395 & T_4329_82;
  assign T_45397 = T_45396 & T_4329_81;
  assign T_45398 = T_45397 & T_4329_80;
  assign T_45399 = T_45398 & T_4329_79;
  assign T_45401 = T_27872 & T_4334_109;
  assign T_45402 = T_45401 & T_4334_108;
  assign T_45403 = T_45402 & T_4334_107;
  assign T_45404 = T_45403 & T_4334_106;
  assign T_45405 = T_45404 & T_4334_105;
  assign T_45406 = T_45405 & T_4334_104;
  assign T_45407 = T_45406 & T_4334_103;
  assign T_45408 = T_45407 & T_4334_102;
  assign T_45409 = T_45408 & T_4334_101;
  assign T_45410 = T_45409 & T_4334_100;
  assign T_45411 = T_45410 & T_4334_99;
  assign T_45412 = T_45411 & T_4334_98;
  assign T_45413 = T_45412 & T_4334_97;
  assign T_45414 = T_45413 & T_4334_96;
  assign T_45415 = T_45414 & T_4334_95;
  assign T_45416 = T_45415 & T_4334_94;
  assign T_45417 = T_45416 & T_4334_93;
  assign T_45418 = T_45417 & T_4334_92;
  assign T_45419 = T_45418 & T_4334_91;
  assign T_45420 = T_45419 & T_4334_90;
  assign T_45421 = T_45420 & T_4334_89;
  assign T_45422 = T_45421 & T_4334_88;
  assign T_45423 = T_45422 & T_4334_87;
  assign T_45424 = T_45423 & T_4334_86;
  assign T_45425 = T_45424 & T_4334_85;
  assign T_45426 = T_45425 & T_4334_84;
  assign T_45427 = T_45426 & T_4334_83;
  assign T_45428 = T_45427 & T_4334_82;
  assign T_45429 = T_45428 & T_4334_81;
  assign T_45430 = T_45429 & T_4334_80;
  assign T_45431 = T_45430 & T_4334_79;
  assign T_45473 = T_26596 & T_4319_140;
  assign T_45474 = T_45473 & T_4319_139;
  assign T_45475 = T_45474 & T_4319_138;
  assign T_45476 = T_45475 & T_4319_137;
  assign T_45477 = T_45476 & T_4319_136;
  assign T_45478 = T_45477 & T_4319_135;
  assign T_45479 = T_45478 & T_4319_134;
  assign T_45480 = T_45479 & T_4319_133;
  assign T_45481 = T_45480 & T_4319_132;
  assign T_45482 = T_45481 & T_4319_131;
  assign T_45483 = T_45482 & T_4319_130;
  assign T_45484 = T_45483 & T_4319_129;
  assign T_45485 = T_45484 & T_4319_128;
  assign T_45486 = T_45485 & T_4319_127;
  assign T_45487 = T_45486 & T_4319_126;
  assign T_45488 = T_45487 & T_4319_125;
  assign T_45489 = T_45488 & T_4319_124;
  assign T_45490 = T_45489 & T_4319_123;
  assign T_45491 = T_45490 & T_4319_122;
  assign T_45493 = T_26602 & T_4324_140;
  assign T_45494 = T_45493 & T_4324_139;
  assign T_45495 = T_45494 & T_4324_138;
  assign T_45496 = T_45495 & T_4324_137;
  assign T_45497 = T_45496 & T_4324_136;
  assign T_45498 = T_45497 & T_4324_135;
  assign T_45499 = T_45498 & T_4324_134;
  assign T_45500 = T_45499 & T_4324_133;
  assign T_45501 = T_45500 & T_4324_132;
  assign T_45502 = T_45501 & T_4324_131;
  assign T_45503 = T_45502 & T_4324_130;
  assign T_45504 = T_45503 & T_4324_129;
  assign T_45505 = T_45504 & T_4324_128;
  assign T_45506 = T_45505 & T_4324_127;
  assign T_45507 = T_45506 & T_4324_126;
  assign T_45508 = T_45507 & T_4324_125;
  assign T_45509 = T_45508 & T_4324_124;
  assign T_45510 = T_45509 & T_4324_123;
  assign T_45511 = T_45510 & T_4324_122;
  assign T_45513 = T_26606 & T_4329_140;
  assign T_45514 = T_45513 & T_4329_139;
  assign T_45515 = T_45514 & T_4329_138;
  assign T_45516 = T_45515 & T_4329_137;
  assign T_45517 = T_45516 & T_4329_136;
  assign T_45518 = T_45517 & T_4329_135;
  assign T_45519 = T_45518 & T_4329_134;
  assign T_45520 = T_45519 & T_4329_133;
  assign T_45521 = T_45520 & T_4329_132;
  assign T_45522 = T_45521 & T_4329_131;
  assign T_45523 = T_45522 & T_4329_130;
  assign T_45524 = T_45523 & T_4329_129;
  assign T_45525 = T_45524 & T_4329_128;
  assign T_45526 = T_45525 & T_4329_127;
  assign T_45527 = T_45526 & T_4329_126;
  assign T_45528 = T_45527 & T_4329_125;
  assign T_45529 = T_45528 & T_4329_124;
  assign T_45530 = T_45529 & T_4329_123;
  assign T_45531 = T_45530 & T_4329_122;
  assign T_45533 = T_26612 & T_4334_140;
  assign T_45534 = T_45533 & T_4334_139;
  assign T_45535 = T_45534 & T_4334_138;
  assign T_45536 = T_45535 & T_4334_137;
  assign T_45537 = T_45536 & T_4334_136;
  assign T_45538 = T_45537 & T_4334_135;
  assign T_45539 = T_45538 & T_4334_134;
  assign T_45540 = T_45539 & T_4334_133;
  assign T_45541 = T_45540 & T_4334_132;
  assign T_45542 = T_45541 & T_4334_131;
  assign T_45543 = T_45542 & T_4334_130;
  assign T_45544 = T_45543 & T_4334_129;
  assign T_45545 = T_45544 & T_4334_128;
  assign T_45546 = T_45545 & T_4334_127;
  assign T_45547 = T_45546 & T_4334_126;
  assign T_45548 = T_45547 & T_4334_125;
  assign T_45549 = T_45548 & T_4334_124;
  assign T_45550 = T_45549 & T_4334_123;
  assign T_45551 = T_45550 & T_4334_122;
  assign T_45571 = T_45490 & T_4319_121;
  assign T_45591 = T_45510 & T_4324_121;
  assign T_45611 = T_45530 & T_4329_121;
  assign T_45631 = T_45550 & T_4334_121;
  assign T_45650 = T_45489 & T_4319_122;
  assign T_45651 = T_45650 & T_4319_121;
  assign T_45670 = T_45509 & T_4324_122;
  assign T_45671 = T_45670 & T_4324_121;
  assign T_45690 = T_45529 & T_4329_122;
  assign T_45691 = T_45690 & T_4329_121;
  assign T_45710 = T_45549 & T_4334_122;
  assign T_45711 = T_45710 & T_4334_121;
  assign T_45729 = T_45488 & T_4319_123;
  assign T_45730 = T_45729 & T_4319_122;
  assign T_45731 = T_45730 & T_4319_121;
  assign T_45749 = T_45508 & T_4324_123;
  assign T_45750 = T_45749 & T_4324_122;
  assign T_45751 = T_45750 & T_4324_121;
  assign T_45769 = T_45528 & T_4329_123;
  assign T_45770 = T_45769 & T_4329_122;
  assign T_45771 = T_45770 & T_4329_121;
  assign T_45789 = T_45548 & T_4334_123;
  assign T_45790 = T_45789 & T_4334_122;
  assign T_45791 = T_45790 & T_4334_121;
  assign T_45808 = T_45487 & T_4319_124;
  assign T_45809 = T_45808 & T_4319_123;
  assign T_45810 = T_45809 & T_4319_122;
  assign T_45811 = T_45810 & T_4319_121;
  assign T_45828 = T_45507 & T_4324_124;
  assign T_45829 = T_45828 & T_4324_123;
  assign T_45830 = T_45829 & T_4324_122;
  assign T_45831 = T_45830 & T_4324_121;
  assign T_45848 = T_45527 & T_4329_124;
  assign T_45849 = T_45848 & T_4329_123;
  assign T_45850 = T_45849 & T_4329_122;
  assign T_45851 = T_45850 & T_4329_121;
  assign T_45868 = T_45547 & T_4334_124;
  assign T_45869 = T_45868 & T_4334_123;
  assign T_45870 = T_45869 & T_4334_122;
  assign T_45871 = T_45870 & T_4334_121;
  assign T_45887 = T_45486 & T_4319_125;
  assign T_45888 = T_45887 & T_4319_124;
  assign T_45889 = T_45888 & T_4319_123;
  assign T_45890 = T_45889 & T_4319_122;
  assign T_45891 = T_45890 & T_4319_121;
  assign T_45907 = T_45506 & T_4324_125;
  assign T_45908 = T_45907 & T_4324_124;
  assign T_45909 = T_45908 & T_4324_123;
  assign T_45910 = T_45909 & T_4324_122;
  assign T_45911 = T_45910 & T_4324_121;
  assign T_45927 = T_45526 & T_4329_125;
  assign T_45928 = T_45927 & T_4329_124;
  assign T_45929 = T_45928 & T_4329_123;
  assign T_45930 = T_45929 & T_4329_122;
  assign T_45931 = T_45930 & T_4329_121;
  assign T_45947 = T_45546 & T_4334_125;
  assign T_45948 = T_45947 & T_4334_124;
  assign T_45949 = T_45948 & T_4334_123;
  assign T_45950 = T_45949 & T_4334_122;
  assign T_45951 = T_45950 & T_4334_121;
  assign T_45966 = T_45485 & T_4319_126;
  assign T_45967 = T_45966 & T_4319_125;
  assign T_45968 = T_45967 & T_4319_124;
  assign T_45969 = T_45968 & T_4319_123;
  assign T_45970 = T_45969 & T_4319_122;
  assign T_45971 = T_45970 & T_4319_121;
  assign T_45986 = T_45505 & T_4324_126;
  assign T_45987 = T_45986 & T_4324_125;
  assign T_45988 = T_45987 & T_4324_124;
  assign T_45989 = T_45988 & T_4324_123;
  assign T_45990 = T_45989 & T_4324_122;
  assign T_45991 = T_45990 & T_4324_121;
  assign T_46006 = T_45525 & T_4329_126;
  assign T_46007 = T_46006 & T_4329_125;
  assign T_46008 = T_46007 & T_4329_124;
  assign T_46009 = T_46008 & T_4329_123;
  assign T_46010 = T_46009 & T_4329_122;
  assign T_46011 = T_46010 & T_4329_121;
  assign T_46026 = T_45545 & T_4334_126;
  assign T_46027 = T_46026 & T_4334_125;
  assign T_46028 = T_46027 & T_4334_124;
  assign T_46029 = T_46028 & T_4334_123;
  assign T_46030 = T_46029 & T_4334_122;
  assign T_46031 = T_46030 & T_4334_121;
  assign T_46045 = T_45484 & T_4319_127;
  assign T_46046 = T_46045 & T_4319_126;
  assign T_46047 = T_46046 & T_4319_125;
  assign T_46048 = T_46047 & T_4319_124;
  assign T_46049 = T_46048 & T_4319_123;
  assign T_46050 = T_46049 & T_4319_122;
  assign T_46051 = T_46050 & T_4319_121;
  assign T_46065 = T_45504 & T_4324_127;
  assign T_46066 = T_46065 & T_4324_126;
  assign T_46067 = T_46066 & T_4324_125;
  assign T_46068 = T_46067 & T_4324_124;
  assign T_46069 = T_46068 & T_4324_123;
  assign T_46070 = T_46069 & T_4324_122;
  assign T_46071 = T_46070 & T_4324_121;
  assign T_46085 = T_45524 & T_4329_127;
  assign T_46086 = T_46085 & T_4329_126;
  assign T_46087 = T_46086 & T_4329_125;
  assign T_46088 = T_46087 & T_4329_124;
  assign T_46089 = T_46088 & T_4329_123;
  assign T_46090 = T_46089 & T_4329_122;
  assign T_46091 = T_46090 & T_4329_121;
  assign T_46105 = T_45544 & T_4334_127;
  assign T_46106 = T_46105 & T_4334_126;
  assign T_46107 = T_46106 & T_4334_125;
  assign T_46108 = T_46107 & T_4334_124;
  assign T_46109 = T_46108 & T_4334_123;
  assign T_46110 = T_46109 & T_4334_122;
  assign T_46111 = T_46110 & T_4334_121;
  assign T_46124 = T_45483 & T_4319_128;
  assign T_46125 = T_46124 & T_4319_127;
  assign T_46126 = T_46125 & T_4319_126;
  assign T_46127 = T_46126 & T_4319_125;
  assign T_46128 = T_46127 & T_4319_124;
  assign T_46129 = T_46128 & T_4319_123;
  assign T_46130 = T_46129 & T_4319_122;
  assign T_46131 = T_46130 & T_4319_121;
  assign T_46144 = T_45503 & T_4324_128;
  assign T_46145 = T_46144 & T_4324_127;
  assign T_46146 = T_46145 & T_4324_126;
  assign T_46147 = T_46146 & T_4324_125;
  assign T_46148 = T_46147 & T_4324_124;
  assign T_46149 = T_46148 & T_4324_123;
  assign T_46150 = T_46149 & T_4324_122;
  assign T_46151 = T_46150 & T_4324_121;
  assign T_46164 = T_45523 & T_4329_128;
  assign T_46165 = T_46164 & T_4329_127;
  assign T_46166 = T_46165 & T_4329_126;
  assign T_46167 = T_46166 & T_4329_125;
  assign T_46168 = T_46167 & T_4329_124;
  assign T_46169 = T_46168 & T_4329_123;
  assign T_46170 = T_46169 & T_4329_122;
  assign T_46171 = T_46170 & T_4329_121;
  assign T_46184 = T_45543 & T_4334_128;
  assign T_46185 = T_46184 & T_4334_127;
  assign T_46186 = T_46185 & T_4334_126;
  assign T_46187 = T_46186 & T_4334_125;
  assign T_46188 = T_46187 & T_4334_124;
  assign T_46189 = T_46188 & T_4334_123;
  assign T_46190 = T_46189 & T_4334_122;
  assign T_46191 = T_46190 & T_4334_121;
  assign T_46203 = T_45482 & T_4319_129;
  assign T_46204 = T_46203 & T_4319_128;
  assign T_46205 = T_46204 & T_4319_127;
  assign T_46206 = T_46205 & T_4319_126;
  assign T_46207 = T_46206 & T_4319_125;
  assign T_46208 = T_46207 & T_4319_124;
  assign T_46209 = T_46208 & T_4319_123;
  assign T_46210 = T_46209 & T_4319_122;
  assign T_46211 = T_46210 & T_4319_121;
  assign T_46223 = T_45502 & T_4324_129;
  assign T_46224 = T_46223 & T_4324_128;
  assign T_46225 = T_46224 & T_4324_127;
  assign T_46226 = T_46225 & T_4324_126;
  assign T_46227 = T_46226 & T_4324_125;
  assign T_46228 = T_46227 & T_4324_124;
  assign T_46229 = T_46228 & T_4324_123;
  assign T_46230 = T_46229 & T_4324_122;
  assign T_46231 = T_46230 & T_4324_121;
  assign T_46243 = T_45522 & T_4329_129;
  assign T_46244 = T_46243 & T_4329_128;
  assign T_46245 = T_46244 & T_4329_127;
  assign T_46246 = T_46245 & T_4329_126;
  assign T_46247 = T_46246 & T_4329_125;
  assign T_46248 = T_46247 & T_4329_124;
  assign T_46249 = T_46248 & T_4329_123;
  assign T_46250 = T_46249 & T_4329_122;
  assign T_46251 = T_46250 & T_4329_121;
  assign T_46263 = T_45542 & T_4334_129;
  assign T_46264 = T_46263 & T_4334_128;
  assign T_46265 = T_46264 & T_4334_127;
  assign T_46266 = T_46265 & T_4334_126;
  assign T_46267 = T_46266 & T_4334_125;
  assign T_46268 = T_46267 & T_4334_124;
  assign T_46269 = T_46268 & T_4334_123;
  assign T_46270 = T_46269 & T_4334_122;
  assign T_46271 = T_46270 & T_4334_121;
  assign T_46282 = T_45481 & T_4319_130;
  assign T_46283 = T_46282 & T_4319_129;
  assign T_46284 = T_46283 & T_4319_128;
  assign T_46285 = T_46284 & T_4319_127;
  assign T_46286 = T_46285 & T_4319_126;
  assign T_46287 = T_46286 & T_4319_125;
  assign T_46288 = T_46287 & T_4319_124;
  assign T_46289 = T_46288 & T_4319_123;
  assign T_46290 = T_46289 & T_4319_122;
  assign T_46291 = T_46290 & T_4319_121;
  assign T_46302 = T_45501 & T_4324_130;
  assign T_46303 = T_46302 & T_4324_129;
  assign T_46304 = T_46303 & T_4324_128;
  assign T_46305 = T_46304 & T_4324_127;
  assign T_46306 = T_46305 & T_4324_126;
  assign T_46307 = T_46306 & T_4324_125;
  assign T_46308 = T_46307 & T_4324_124;
  assign T_46309 = T_46308 & T_4324_123;
  assign T_46310 = T_46309 & T_4324_122;
  assign T_46311 = T_46310 & T_4324_121;
  assign T_46322 = T_45521 & T_4329_130;
  assign T_46323 = T_46322 & T_4329_129;
  assign T_46324 = T_46323 & T_4329_128;
  assign T_46325 = T_46324 & T_4329_127;
  assign T_46326 = T_46325 & T_4329_126;
  assign T_46327 = T_46326 & T_4329_125;
  assign T_46328 = T_46327 & T_4329_124;
  assign T_46329 = T_46328 & T_4329_123;
  assign T_46330 = T_46329 & T_4329_122;
  assign T_46331 = T_46330 & T_4329_121;
  assign T_46342 = T_45541 & T_4334_130;
  assign T_46343 = T_46342 & T_4334_129;
  assign T_46344 = T_46343 & T_4334_128;
  assign T_46345 = T_46344 & T_4334_127;
  assign T_46346 = T_46345 & T_4334_126;
  assign T_46347 = T_46346 & T_4334_125;
  assign T_46348 = T_46347 & T_4334_124;
  assign T_46349 = T_46348 & T_4334_123;
  assign T_46350 = T_46349 & T_4334_122;
  assign T_46351 = T_46350 & T_4334_121;
  assign T_46361 = T_45480 & T_4319_131;
  assign T_46362 = T_46361 & T_4319_130;
  assign T_46363 = T_46362 & T_4319_129;
  assign T_46364 = T_46363 & T_4319_128;
  assign T_46365 = T_46364 & T_4319_127;
  assign T_46366 = T_46365 & T_4319_126;
  assign T_46367 = T_46366 & T_4319_125;
  assign T_46368 = T_46367 & T_4319_124;
  assign T_46369 = T_46368 & T_4319_123;
  assign T_46370 = T_46369 & T_4319_122;
  assign T_46371 = T_46370 & T_4319_121;
  assign T_46381 = T_45500 & T_4324_131;
  assign T_46382 = T_46381 & T_4324_130;
  assign T_46383 = T_46382 & T_4324_129;
  assign T_46384 = T_46383 & T_4324_128;
  assign T_46385 = T_46384 & T_4324_127;
  assign T_46386 = T_46385 & T_4324_126;
  assign T_46387 = T_46386 & T_4324_125;
  assign T_46388 = T_46387 & T_4324_124;
  assign T_46389 = T_46388 & T_4324_123;
  assign T_46390 = T_46389 & T_4324_122;
  assign T_46391 = T_46390 & T_4324_121;
  assign T_46401 = T_45520 & T_4329_131;
  assign T_46402 = T_46401 & T_4329_130;
  assign T_46403 = T_46402 & T_4329_129;
  assign T_46404 = T_46403 & T_4329_128;
  assign T_46405 = T_46404 & T_4329_127;
  assign T_46406 = T_46405 & T_4329_126;
  assign T_46407 = T_46406 & T_4329_125;
  assign T_46408 = T_46407 & T_4329_124;
  assign T_46409 = T_46408 & T_4329_123;
  assign T_46410 = T_46409 & T_4329_122;
  assign T_46411 = T_46410 & T_4329_121;
  assign T_46421 = T_45540 & T_4334_131;
  assign T_46422 = T_46421 & T_4334_130;
  assign T_46423 = T_46422 & T_4334_129;
  assign T_46424 = T_46423 & T_4334_128;
  assign T_46425 = T_46424 & T_4334_127;
  assign T_46426 = T_46425 & T_4334_126;
  assign T_46427 = T_46426 & T_4334_125;
  assign T_46428 = T_46427 & T_4334_124;
  assign T_46429 = T_46428 & T_4334_123;
  assign T_46430 = T_46429 & T_4334_122;
  assign T_46431 = T_46430 & T_4334_121;
  assign T_46440 = T_45479 & T_4319_132;
  assign T_46441 = T_46440 & T_4319_131;
  assign T_46442 = T_46441 & T_4319_130;
  assign T_46443 = T_46442 & T_4319_129;
  assign T_46444 = T_46443 & T_4319_128;
  assign T_46445 = T_46444 & T_4319_127;
  assign T_46446 = T_46445 & T_4319_126;
  assign T_46447 = T_46446 & T_4319_125;
  assign T_46448 = T_46447 & T_4319_124;
  assign T_46449 = T_46448 & T_4319_123;
  assign T_46450 = T_46449 & T_4319_122;
  assign T_46451 = T_46450 & T_4319_121;
  assign T_46460 = T_45499 & T_4324_132;
  assign T_46461 = T_46460 & T_4324_131;
  assign T_46462 = T_46461 & T_4324_130;
  assign T_46463 = T_46462 & T_4324_129;
  assign T_46464 = T_46463 & T_4324_128;
  assign T_46465 = T_46464 & T_4324_127;
  assign T_46466 = T_46465 & T_4324_126;
  assign T_46467 = T_46466 & T_4324_125;
  assign T_46468 = T_46467 & T_4324_124;
  assign T_46469 = T_46468 & T_4324_123;
  assign T_46470 = T_46469 & T_4324_122;
  assign T_46471 = T_46470 & T_4324_121;
  assign T_46480 = T_45519 & T_4329_132;
  assign T_46481 = T_46480 & T_4329_131;
  assign T_46482 = T_46481 & T_4329_130;
  assign T_46483 = T_46482 & T_4329_129;
  assign T_46484 = T_46483 & T_4329_128;
  assign T_46485 = T_46484 & T_4329_127;
  assign T_46486 = T_46485 & T_4329_126;
  assign T_46487 = T_46486 & T_4329_125;
  assign T_46488 = T_46487 & T_4329_124;
  assign T_46489 = T_46488 & T_4329_123;
  assign T_46490 = T_46489 & T_4329_122;
  assign T_46491 = T_46490 & T_4329_121;
  assign T_46500 = T_45539 & T_4334_132;
  assign T_46501 = T_46500 & T_4334_131;
  assign T_46502 = T_46501 & T_4334_130;
  assign T_46503 = T_46502 & T_4334_129;
  assign T_46504 = T_46503 & T_4334_128;
  assign T_46505 = T_46504 & T_4334_127;
  assign T_46506 = T_46505 & T_4334_126;
  assign T_46507 = T_46506 & T_4334_125;
  assign T_46508 = T_46507 & T_4334_124;
  assign T_46509 = T_46508 & T_4334_123;
  assign T_46510 = T_46509 & T_4334_122;
  assign T_46511 = T_46510 & T_4334_121;
  assign T_46519 = T_45478 & T_4319_133;
  assign T_46520 = T_46519 & T_4319_132;
  assign T_46521 = T_46520 & T_4319_131;
  assign T_46522 = T_46521 & T_4319_130;
  assign T_46523 = T_46522 & T_4319_129;
  assign T_46524 = T_46523 & T_4319_128;
  assign T_46525 = T_46524 & T_4319_127;
  assign T_46526 = T_46525 & T_4319_126;
  assign T_46527 = T_46526 & T_4319_125;
  assign T_46528 = T_46527 & T_4319_124;
  assign T_46529 = T_46528 & T_4319_123;
  assign T_46530 = T_46529 & T_4319_122;
  assign T_46531 = T_46530 & T_4319_121;
  assign T_46539 = T_45498 & T_4324_133;
  assign T_46540 = T_46539 & T_4324_132;
  assign T_46541 = T_46540 & T_4324_131;
  assign T_46542 = T_46541 & T_4324_130;
  assign T_46543 = T_46542 & T_4324_129;
  assign T_46544 = T_46543 & T_4324_128;
  assign T_46545 = T_46544 & T_4324_127;
  assign T_46546 = T_46545 & T_4324_126;
  assign T_46547 = T_46546 & T_4324_125;
  assign T_46548 = T_46547 & T_4324_124;
  assign T_46549 = T_46548 & T_4324_123;
  assign T_46550 = T_46549 & T_4324_122;
  assign T_46551 = T_46550 & T_4324_121;
  assign T_46559 = T_45518 & T_4329_133;
  assign T_46560 = T_46559 & T_4329_132;
  assign T_46561 = T_46560 & T_4329_131;
  assign T_46562 = T_46561 & T_4329_130;
  assign T_46563 = T_46562 & T_4329_129;
  assign T_46564 = T_46563 & T_4329_128;
  assign T_46565 = T_46564 & T_4329_127;
  assign T_46566 = T_46565 & T_4329_126;
  assign T_46567 = T_46566 & T_4329_125;
  assign T_46568 = T_46567 & T_4329_124;
  assign T_46569 = T_46568 & T_4329_123;
  assign T_46570 = T_46569 & T_4329_122;
  assign T_46571 = T_46570 & T_4329_121;
  assign T_46579 = T_45538 & T_4334_133;
  assign T_46580 = T_46579 & T_4334_132;
  assign T_46581 = T_46580 & T_4334_131;
  assign T_46582 = T_46581 & T_4334_130;
  assign T_46583 = T_46582 & T_4334_129;
  assign T_46584 = T_46583 & T_4334_128;
  assign T_46585 = T_46584 & T_4334_127;
  assign T_46586 = T_46585 & T_4334_126;
  assign T_46587 = T_46586 & T_4334_125;
  assign T_46588 = T_46587 & T_4334_124;
  assign T_46589 = T_46588 & T_4334_123;
  assign T_46590 = T_46589 & T_4334_122;
  assign T_46591 = T_46590 & T_4334_121;
  assign T_46598 = T_45477 & T_4319_134;
  assign T_46599 = T_46598 & T_4319_133;
  assign T_46600 = T_46599 & T_4319_132;
  assign T_46601 = T_46600 & T_4319_131;
  assign T_46602 = T_46601 & T_4319_130;
  assign T_46603 = T_46602 & T_4319_129;
  assign T_46604 = T_46603 & T_4319_128;
  assign T_46605 = T_46604 & T_4319_127;
  assign T_46606 = T_46605 & T_4319_126;
  assign T_46607 = T_46606 & T_4319_125;
  assign T_46608 = T_46607 & T_4319_124;
  assign T_46609 = T_46608 & T_4319_123;
  assign T_46610 = T_46609 & T_4319_122;
  assign T_46611 = T_46610 & T_4319_121;
  assign T_46618 = T_45497 & T_4324_134;
  assign T_46619 = T_46618 & T_4324_133;
  assign T_46620 = T_46619 & T_4324_132;
  assign T_46621 = T_46620 & T_4324_131;
  assign T_46622 = T_46621 & T_4324_130;
  assign T_46623 = T_46622 & T_4324_129;
  assign T_46624 = T_46623 & T_4324_128;
  assign T_46625 = T_46624 & T_4324_127;
  assign T_46626 = T_46625 & T_4324_126;
  assign T_46627 = T_46626 & T_4324_125;
  assign T_46628 = T_46627 & T_4324_124;
  assign T_46629 = T_46628 & T_4324_123;
  assign T_46630 = T_46629 & T_4324_122;
  assign T_46631 = T_46630 & T_4324_121;
  assign T_46638 = T_45517 & T_4329_134;
  assign T_46639 = T_46638 & T_4329_133;
  assign T_46640 = T_46639 & T_4329_132;
  assign T_46641 = T_46640 & T_4329_131;
  assign T_46642 = T_46641 & T_4329_130;
  assign T_46643 = T_46642 & T_4329_129;
  assign T_46644 = T_46643 & T_4329_128;
  assign T_46645 = T_46644 & T_4329_127;
  assign T_46646 = T_46645 & T_4329_126;
  assign T_46647 = T_46646 & T_4329_125;
  assign T_46648 = T_46647 & T_4329_124;
  assign T_46649 = T_46648 & T_4329_123;
  assign T_46650 = T_46649 & T_4329_122;
  assign T_46651 = T_46650 & T_4329_121;
  assign T_46658 = T_45537 & T_4334_134;
  assign T_46659 = T_46658 & T_4334_133;
  assign T_46660 = T_46659 & T_4334_132;
  assign T_46661 = T_46660 & T_4334_131;
  assign T_46662 = T_46661 & T_4334_130;
  assign T_46663 = T_46662 & T_4334_129;
  assign T_46664 = T_46663 & T_4334_128;
  assign T_46665 = T_46664 & T_4334_127;
  assign T_46666 = T_46665 & T_4334_126;
  assign T_46667 = T_46666 & T_4334_125;
  assign T_46668 = T_46667 & T_4334_124;
  assign T_46669 = T_46668 & T_4334_123;
  assign T_46670 = T_46669 & T_4334_122;
  assign T_46671 = T_46670 & T_4334_121;
  assign T_46677 = T_45476 & T_4319_135;
  assign T_46678 = T_46677 & T_4319_134;
  assign T_46679 = T_46678 & T_4319_133;
  assign T_46680 = T_46679 & T_4319_132;
  assign T_46681 = T_46680 & T_4319_131;
  assign T_46682 = T_46681 & T_4319_130;
  assign T_46683 = T_46682 & T_4319_129;
  assign T_46684 = T_46683 & T_4319_128;
  assign T_46685 = T_46684 & T_4319_127;
  assign T_46686 = T_46685 & T_4319_126;
  assign T_46687 = T_46686 & T_4319_125;
  assign T_46688 = T_46687 & T_4319_124;
  assign T_46689 = T_46688 & T_4319_123;
  assign T_46690 = T_46689 & T_4319_122;
  assign T_46691 = T_46690 & T_4319_121;
  assign T_46697 = T_45496 & T_4324_135;
  assign T_46698 = T_46697 & T_4324_134;
  assign T_46699 = T_46698 & T_4324_133;
  assign T_46700 = T_46699 & T_4324_132;
  assign T_46701 = T_46700 & T_4324_131;
  assign T_46702 = T_46701 & T_4324_130;
  assign T_46703 = T_46702 & T_4324_129;
  assign T_46704 = T_46703 & T_4324_128;
  assign T_46705 = T_46704 & T_4324_127;
  assign T_46706 = T_46705 & T_4324_126;
  assign T_46707 = T_46706 & T_4324_125;
  assign T_46708 = T_46707 & T_4324_124;
  assign T_46709 = T_46708 & T_4324_123;
  assign T_46710 = T_46709 & T_4324_122;
  assign T_46711 = T_46710 & T_4324_121;
  assign T_46717 = T_45516 & T_4329_135;
  assign T_46718 = T_46717 & T_4329_134;
  assign T_46719 = T_46718 & T_4329_133;
  assign T_46720 = T_46719 & T_4329_132;
  assign T_46721 = T_46720 & T_4329_131;
  assign T_46722 = T_46721 & T_4329_130;
  assign T_46723 = T_46722 & T_4329_129;
  assign T_46724 = T_46723 & T_4329_128;
  assign T_46725 = T_46724 & T_4329_127;
  assign T_46726 = T_46725 & T_4329_126;
  assign T_46727 = T_46726 & T_4329_125;
  assign T_46728 = T_46727 & T_4329_124;
  assign T_46729 = T_46728 & T_4329_123;
  assign T_46730 = T_46729 & T_4329_122;
  assign T_46731 = T_46730 & T_4329_121;
  assign T_46737 = T_45536 & T_4334_135;
  assign T_46738 = T_46737 & T_4334_134;
  assign T_46739 = T_46738 & T_4334_133;
  assign T_46740 = T_46739 & T_4334_132;
  assign T_46741 = T_46740 & T_4334_131;
  assign T_46742 = T_46741 & T_4334_130;
  assign T_46743 = T_46742 & T_4334_129;
  assign T_46744 = T_46743 & T_4334_128;
  assign T_46745 = T_46744 & T_4334_127;
  assign T_46746 = T_46745 & T_4334_126;
  assign T_46747 = T_46746 & T_4334_125;
  assign T_46748 = T_46747 & T_4334_124;
  assign T_46749 = T_46748 & T_4334_123;
  assign T_46750 = T_46749 & T_4334_122;
  assign T_46751 = T_46750 & T_4334_121;
  assign T_46756 = T_45475 & T_4319_136;
  assign T_46757 = T_46756 & T_4319_135;
  assign T_46758 = T_46757 & T_4319_134;
  assign T_46759 = T_46758 & T_4319_133;
  assign T_46760 = T_46759 & T_4319_132;
  assign T_46761 = T_46760 & T_4319_131;
  assign T_46762 = T_46761 & T_4319_130;
  assign T_46763 = T_46762 & T_4319_129;
  assign T_46764 = T_46763 & T_4319_128;
  assign T_46765 = T_46764 & T_4319_127;
  assign T_46766 = T_46765 & T_4319_126;
  assign T_46767 = T_46766 & T_4319_125;
  assign T_46768 = T_46767 & T_4319_124;
  assign T_46769 = T_46768 & T_4319_123;
  assign T_46770 = T_46769 & T_4319_122;
  assign T_46771 = T_46770 & T_4319_121;
  assign T_46776 = T_45495 & T_4324_136;
  assign T_46777 = T_46776 & T_4324_135;
  assign T_46778 = T_46777 & T_4324_134;
  assign T_46779 = T_46778 & T_4324_133;
  assign T_46780 = T_46779 & T_4324_132;
  assign T_46781 = T_46780 & T_4324_131;
  assign T_46782 = T_46781 & T_4324_130;
  assign T_46783 = T_46782 & T_4324_129;
  assign T_46784 = T_46783 & T_4324_128;
  assign T_46785 = T_46784 & T_4324_127;
  assign T_46786 = T_46785 & T_4324_126;
  assign T_46787 = T_46786 & T_4324_125;
  assign T_46788 = T_46787 & T_4324_124;
  assign T_46789 = T_46788 & T_4324_123;
  assign T_46790 = T_46789 & T_4324_122;
  assign T_46791 = T_46790 & T_4324_121;
  assign T_46796 = T_45515 & T_4329_136;
  assign T_46797 = T_46796 & T_4329_135;
  assign T_46798 = T_46797 & T_4329_134;
  assign T_46799 = T_46798 & T_4329_133;
  assign T_46800 = T_46799 & T_4329_132;
  assign T_46801 = T_46800 & T_4329_131;
  assign T_46802 = T_46801 & T_4329_130;
  assign T_46803 = T_46802 & T_4329_129;
  assign T_46804 = T_46803 & T_4329_128;
  assign T_46805 = T_46804 & T_4329_127;
  assign T_46806 = T_46805 & T_4329_126;
  assign T_46807 = T_46806 & T_4329_125;
  assign T_46808 = T_46807 & T_4329_124;
  assign T_46809 = T_46808 & T_4329_123;
  assign T_46810 = T_46809 & T_4329_122;
  assign T_46811 = T_46810 & T_4329_121;
  assign T_46816 = T_45535 & T_4334_136;
  assign T_46817 = T_46816 & T_4334_135;
  assign T_46818 = T_46817 & T_4334_134;
  assign T_46819 = T_46818 & T_4334_133;
  assign T_46820 = T_46819 & T_4334_132;
  assign T_46821 = T_46820 & T_4334_131;
  assign T_46822 = T_46821 & T_4334_130;
  assign T_46823 = T_46822 & T_4334_129;
  assign T_46824 = T_46823 & T_4334_128;
  assign T_46825 = T_46824 & T_4334_127;
  assign T_46826 = T_46825 & T_4334_126;
  assign T_46827 = T_46826 & T_4334_125;
  assign T_46828 = T_46827 & T_4334_124;
  assign T_46829 = T_46828 & T_4334_123;
  assign T_46830 = T_46829 & T_4334_122;
  assign T_46831 = T_46830 & T_4334_121;
  assign T_46835 = T_45474 & T_4319_137;
  assign T_46836 = T_46835 & T_4319_136;
  assign T_46837 = T_46836 & T_4319_135;
  assign T_46838 = T_46837 & T_4319_134;
  assign T_46839 = T_46838 & T_4319_133;
  assign T_46840 = T_46839 & T_4319_132;
  assign T_46841 = T_46840 & T_4319_131;
  assign T_46842 = T_46841 & T_4319_130;
  assign T_46843 = T_46842 & T_4319_129;
  assign T_46844 = T_46843 & T_4319_128;
  assign T_46845 = T_46844 & T_4319_127;
  assign T_46846 = T_46845 & T_4319_126;
  assign T_46847 = T_46846 & T_4319_125;
  assign T_46848 = T_46847 & T_4319_124;
  assign T_46849 = T_46848 & T_4319_123;
  assign T_46850 = T_46849 & T_4319_122;
  assign T_46851 = T_46850 & T_4319_121;
  assign T_46855 = T_45494 & T_4324_137;
  assign T_46856 = T_46855 & T_4324_136;
  assign T_46857 = T_46856 & T_4324_135;
  assign T_46858 = T_46857 & T_4324_134;
  assign T_46859 = T_46858 & T_4324_133;
  assign T_46860 = T_46859 & T_4324_132;
  assign T_46861 = T_46860 & T_4324_131;
  assign T_46862 = T_46861 & T_4324_130;
  assign T_46863 = T_46862 & T_4324_129;
  assign T_46864 = T_46863 & T_4324_128;
  assign T_46865 = T_46864 & T_4324_127;
  assign T_46866 = T_46865 & T_4324_126;
  assign T_46867 = T_46866 & T_4324_125;
  assign T_46868 = T_46867 & T_4324_124;
  assign T_46869 = T_46868 & T_4324_123;
  assign T_46870 = T_46869 & T_4324_122;
  assign T_46871 = T_46870 & T_4324_121;
  assign T_46875 = T_45514 & T_4329_137;
  assign T_46876 = T_46875 & T_4329_136;
  assign T_46877 = T_46876 & T_4329_135;
  assign T_46878 = T_46877 & T_4329_134;
  assign T_46879 = T_46878 & T_4329_133;
  assign T_46880 = T_46879 & T_4329_132;
  assign T_46881 = T_46880 & T_4329_131;
  assign T_46882 = T_46881 & T_4329_130;
  assign T_46883 = T_46882 & T_4329_129;
  assign T_46884 = T_46883 & T_4329_128;
  assign T_46885 = T_46884 & T_4329_127;
  assign T_46886 = T_46885 & T_4329_126;
  assign T_46887 = T_46886 & T_4329_125;
  assign T_46888 = T_46887 & T_4329_124;
  assign T_46889 = T_46888 & T_4329_123;
  assign T_46890 = T_46889 & T_4329_122;
  assign T_46891 = T_46890 & T_4329_121;
  assign T_46895 = T_45534 & T_4334_137;
  assign T_46896 = T_46895 & T_4334_136;
  assign T_46897 = T_46896 & T_4334_135;
  assign T_46898 = T_46897 & T_4334_134;
  assign T_46899 = T_46898 & T_4334_133;
  assign T_46900 = T_46899 & T_4334_132;
  assign T_46901 = T_46900 & T_4334_131;
  assign T_46902 = T_46901 & T_4334_130;
  assign T_46903 = T_46902 & T_4334_129;
  assign T_46904 = T_46903 & T_4334_128;
  assign T_46905 = T_46904 & T_4334_127;
  assign T_46906 = T_46905 & T_4334_126;
  assign T_46907 = T_46906 & T_4334_125;
  assign T_46908 = T_46907 & T_4334_124;
  assign T_46909 = T_46908 & T_4334_123;
  assign T_46910 = T_46909 & T_4334_122;
  assign T_46911 = T_46910 & T_4334_121;
  assign T_46914 = T_45473 & T_4319_138;
  assign T_46915 = T_46914 & T_4319_137;
  assign T_46916 = T_46915 & T_4319_136;
  assign T_46917 = T_46916 & T_4319_135;
  assign T_46918 = T_46917 & T_4319_134;
  assign T_46919 = T_46918 & T_4319_133;
  assign T_46920 = T_46919 & T_4319_132;
  assign T_46921 = T_46920 & T_4319_131;
  assign T_46922 = T_46921 & T_4319_130;
  assign T_46923 = T_46922 & T_4319_129;
  assign T_46924 = T_46923 & T_4319_128;
  assign T_46925 = T_46924 & T_4319_127;
  assign T_46926 = T_46925 & T_4319_126;
  assign T_46927 = T_46926 & T_4319_125;
  assign T_46928 = T_46927 & T_4319_124;
  assign T_46929 = T_46928 & T_4319_123;
  assign T_46930 = T_46929 & T_4319_122;
  assign T_46931 = T_46930 & T_4319_121;
  assign T_46934 = T_45493 & T_4324_138;
  assign T_46935 = T_46934 & T_4324_137;
  assign T_46936 = T_46935 & T_4324_136;
  assign T_46937 = T_46936 & T_4324_135;
  assign T_46938 = T_46937 & T_4324_134;
  assign T_46939 = T_46938 & T_4324_133;
  assign T_46940 = T_46939 & T_4324_132;
  assign T_46941 = T_46940 & T_4324_131;
  assign T_46942 = T_46941 & T_4324_130;
  assign T_46943 = T_46942 & T_4324_129;
  assign T_46944 = T_46943 & T_4324_128;
  assign T_46945 = T_46944 & T_4324_127;
  assign T_46946 = T_46945 & T_4324_126;
  assign T_46947 = T_46946 & T_4324_125;
  assign T_46948 = T_46947 & T_4324_124;
  assign T_46949 = T_46948 & T_4324_123;
  assign T_46950 = T_46949 & T_4324_122;
  assign T_46951 = T_46950 & T_4324_121;
  assign T_46954 = T_45513 & T_4329_138;
  assign T_46955 = T_46954 & T_4329_137;
  assign T_46956 = T_46955 & T_4329_136;
  assign T_46957 = T_46956 & T_4329_135;
  assign T_46958 = T_46957 & T_4329_134;
  assign T_46959 = T_46958 & T_4329_133;
  assign T_46960 = T_46959 & T_4329_132;
  assign T_46961 = T_46960 & T_4329_131;
  assign T_46962 = T_46961 & T_4329_130;
  assign T_46963 = T_46962 & T_4329_129;
  assign T_46964 = T_46963 & T_4329_128;
  assign T_46965 = T_46964 & T_4329_127;
  assign T_46966 = T_46965 & T_4329_126;
  assign T_46967 = T_46966 & T_4329_125;
  assign T_46968 = T_46967 & T_4329_124;
  assign T_46969 = T_46968 & T_4329_123;
  assign T_46970 = T_46969 & T_4329_122;
  assign T_46971 = T_46970 & T_4329_121;
  assign T_46974 = T_45533 & T_4334_138;
  assign T_46975 = T_46974 & T_4334_137;
  assign T_46976 = T_46975 & T_4334_136;
  assign T_46977 = T_46976 & T_4334_135;
  assign T_46978 = T_46977 & T_4334_134;
  assign T_46979 = T_46978 & T_4334_133;
  assign T_46980 = T_46979 & T_4334_132;
  assign T_46981 = T_46980 & T_4334_131;
  assign T_46982 = T_46981 & T_4334_130;
  assign T_46983 = T_46982 & T_4334_129;
  assign T_46984 = T_46983 & T_4334_128;
  assign T_46985 = T_46984 & T_4334_127;
  assign T_46986 = T_46985 & T_4334_126;
  assign T_46987 = T_46986 & T_4334_125;
  assign T_46988 = T_46987 & T_4334_124;
  assign T_46989 = T_46988 & T_4334_123;
  assign T_46990 = T_46989 & T_4334_122;
  assign T_46991 = T_46990 & T_4334_121;
  assign T_46993 = T_26596 & T_4319_139;
  assign T_46994 = T_46993 & T_4319_138;
  assign T_46995 = T_46994 & T_4319_137;
  assign T_46996 = T_46995 & T_4319_136;
  assign T_46997 = T_46996 & T_4319_135;
  assign T_46998 = T_46997 & T_4319_134;
  assign T_46999 = T_46998 & T_4319_133;
  assign T_47000 = T_46999 & T_4319_132;
  assign T_47001 = T_47000 & T_4319_131;
  assign T_47002 = T_47001 & T_4319_130;
  assign T_47003 = T_47002 & T_4319_129;
  assign T_47004 = T_47003 & T_4319_128;
  assign T_47005 = T_47004 & T_4319_127;
  assign T_47006 = T_47005 & T_4319_126;
  assign T_47007 = T_47006 & T_4319_125;
  assign T_47008 = T_47007 & T_4319_124;
  assign T_47009 = T_47008 & T_4319_123;
  assign T_47010 = T_47009 & T_4319_122;
  assign T_47011 = T_47010 & T_4319_121;
  assign T_47013 = T_26602 & T_4324_139;
  assign T_47014 = T_47013 & T_4324_138;
  assign T_47015 = T_47014 & T_4324_137;
  assign T_47016 = T_47015 & T_4324_136;
  assign T_47017 = T_47016 & T_4324_135;
  assign T_47018 = T_47017 & T_4324_134;
  assign T_47019 = T_47018 & T_4324_133;
  assign T_47020 = T_47019 & T_4324_132;
  assign T_47021 = T_47020 & T_4324_131;
  assign T_47022 = T_47021 & T_4324_130;
  assign T_47023 = T_47022 & T_4324_129;
  assign T_47024 = T_47023 & T_4324_128;
  assign T_47025 = T_47024 & T_4324_127;
  assign T_47026 = T_47025 & T_4324_126;
  assign T_47027 = T_47026 & T_4324_125;
  assign T_47028 = T_47027 & T_4324_124;
  assign T_47029 = T_47028 & T_4324_123;
  assign T_47030 = T_47029 & T_4324_122;
  assign T_47031 = T_47030 & T_4324_121;
  assign T_47033 = T_26606 & T_4329_139;
  assign T_47034 = T_47033 & T_4329_138;
  assign T_47035 = T_47034 & T_4329_137;
  assign T_47036 = T_47035 & T_4329_136;
  assign T_47037 = T_47036 & T_4329_135;
  assign T_47038 = T_47037 & T_4329_134;
  assign T_47039 = T_47038 & T_4329_133;
  assign T_47040 = T_47039 & T_4329_132;
  assign T_47041 = T_47040 & T_4329_131;
  assign T_47042 = T_47041 & T_4329_130;
  assign T_47043 = T_47042 & T_4329_129;
  assign T_47044 = T_47043 & T_4329_128;
  assign T_47045 = T_47044 & T_4329_127;
  assign T_47046 = T_47045 & T_4329_126;
  assign T_47047 = T_47046 & T_4329_125;
  assign T_47048 = T_47047 & T_4329_124;
  assign T_47049 = T_47048 & T_4329_123;
  assign T_47050 = T_47049 & T_4329_122;
  assign T_47051 = T_47050 & T_4329_121;
  assign T_47053 = T_26612 & T_4334_139;
  assign T_47054 = T_47053 & T_4334_138;
  assign T_47055 = T_47054 & T_4334_137;
  assign T_47056 = T_47055 & T_4334_136;
  assign T_47057 = T_47056 & T_4334_135;
  assign T_47058 = T_47057 & T_4334_134;
  assign T_47059 = T_47058 & T_4334_133;
  assign T_47060 = T_47059 & T_4334_132;
  assign T_47061 = T_47060 & T_4334_131;
  assign T_47062 = T_47061 & T_4334_130;
  assign T_47063 = T_47062 & T_4334_129;
  assign T_47064 = T_47063 & T_4334_128;
  assign T_47065 = T_47064 & T_4334_127;
  assign T_47066 = T_47065 & T_4334_126;
  assign T_47067 = T_47066 & T_4334_125;
  assign T_47068 = T_47067 & T_4334_124;
  assign T_47069 = T_47068 & T_4334_123;
  assign T_47070 = T_47069 & T_4334_122;
  assign T_47071 = T_47070 & T_4334_121;
  assign T_47656_0 = 1'h1;
  assign T_47656_1 = 1'h1;
  assign T_47656_2 = 1'h1;
  assign T_47656_3 = 1'h1;
  assign T_47656_4 = 1'h1;
  assign T_47656_5 = 1'h1;
  assign T_47656_6 = 1'h1;
  assign T_47656_7 = 1'h1;
  assign T_47656_8 = 1'h1;
  assign T_47656_9 = 1'h1;
  assign T_47656_10 = 1'h1;
  assign T_47656_11 = 1'h1;
  assign T_47656_12 = 1'h1;
  assign T_47656_13 = 1'h1;
  assign T_47656_14 = 1'h1;
  assign T_47656_15 = 1'h1;
  assign T_47656_16 = 1'h1;
  assign T_47656_17 = 1'h1;
  assign T_47656_18 = 1'h1;
  assign T_47656_19 = 1'h1;
  assign T_47656_20 = 1'h1;
  assign T_47656_21 = 1'h1;
  assign T_47656_22 = 1'h1;
  assign T_47656_23 = 1'h1;
  assign T_47656_24 = 1'h1;
  assign T_47656_25 = 1'h1;
  assign T_47656_26 = 1'h1;
  assign T_47656_27 = 1'h1;
  assign T_47656_28 = 1'h1;
  assign T_47656_29 = 1'h1;
  assign T_47656_30 = 1'h1;
  assign T_47656_31 = 1'h1;
  assign T_47656_32 = 1'h1;
  assign T_47656_33 = 1'h1;
  assign T_47656_34 = 1'h1;
  assign T_47656_35 = 1'h1;
  assign T_47656_36 = 1'h1;
  assign T_47656_37 = 1'h1;
  assign T_47656_38 = 1'h1;
  assign T_47656_39 = 1'h1;
  assign T_47656_40 = 1'h1;
  assign T_47656_41 = 1'h1;
  assign T_47656_42 = 1'h1;
  assign T_47656_43 = 1'h1;
  assign T_47656_44 = 1'h1;
  assign T_47656_45 = 1'h1;
  assign T_47656_46 = 1'h1;
  assign T_47656_47 = 1'h1;
  assign T_47656_48 = 1'h1;
  assign T_47656_49 = 1'h1;
  assign T_47656_50 = 1'h1;
  assign T_47656_51 = 1'h1;
  assign T_47656_52 = 1'h1;
  assign T_47656_53 = 1'h1;
  assign T_47656_54 = 1'h1;
  assign T_47656_55 = 1'h1;
  assign T_47656_56 = 1'h1;
  assign T_47656_57 = 1'h1;
  assign T_47656_58 = 1'h1;
  assign T_47656_59 = 1'h1;
  assign T_47656_60 = 1'h1;
  assign T_47656_61 = 1'h1;
  assign T_47656_62 = 1'h1;
  assign T_47656_63 = 1'h1;
  assign T_47656_64 = 1'h1;
  assign T_47656_65 = 1'h1;
  assign T_47656_66 = 1'h1;
  assign T_47656_67 = 1'h1;
  assign T_47656_68 = 1'h1;
  assign T_47656_69 = 1'h1;
  assign T_47656_70 = 1'h1;
  assign T_47656_71 = 1'h1;
  assign T_47656_72 = 1'h1;
  assign T_47656_73 = 1'h1;
  assign T_47656_74 = 1'h1;
  assign T_47656_75 = 1'h1;
  assign T_47656_76 = 1'h1;
  assign T_47656_77 = 1'h1;
  assign T_47656_78 = 1'h1;
  assign T_47656_79 = 1'h1;
  assign T_47656_80 = 1'h1;
  assign T_47656_81 = 1'h1;
  assign T_47656_82 = 1'h1;
  assign T_47656_83 = 1'h1;
  assign T_47656_84 = 1'h1;
  assign T_47656_85 = 1'h1;
  assign T_47656_86 = 1'h1;
  assign T_47656_87 = 1'h1;
  assign T_47656_88 = 1'h1;
  assign T_47656_89 = 1'h1;
  assign T_47656_90 = 1'h1;
  assign T_47656_91 = 1'h1;
  assign T_47656_92 = 1'h1;
  assign T_47656_93 = 1'h1;
  assign T_47656_94 = 1'h1;
  assign T_47656_95 = 1'h1;
  assign T_47656_96 = 1'h1;
  assign T_47656_97 = 1'h1;
  assign T_47656_98 = 1'h1;
  assign T_47656_99 = 1'h1;
  assign T_47656_100 = 1'h1;
  assign T_47656_101 = 1'h1;
  assign T_47656_102 = 1'h1;
  assign T_47656_103 = 1'h1;
  assign T_47656_104 = 1'h1;
  assign T_47656_105 = 1'h1;
  assign T_47656_106 = 1'h1;
  assign T_47656_107 = 1'h1;
  assign T_47656_108 = 1'h1;
  assign T_47656_109 = 1'h1;
  assign T_47656_110 = 1'h1;
  assign T_47656_111 = 1'h1;
  assign T_47656_112 = 1'h1;
  assign T_47656_113 = 1'h1;
  assign T_47656_114 = 1'h1;
  assign T_47656_115 = 1'h1;
  assign T_47656_116 = 1'h1;
  assign T_47656_117 = 1'h1;
  assign T_47656_118 = 1'h1;
  assign T_47656_119 = 1'h1;
  assign T_47656_120 = 1'h1;
  assign T_47656_121 = 1'h1;
  assign T_47656_122 = 1'h1;
  assign T_47656_123 = 1'h1;
  assign T_47656_124 = 1'h1;
  assign T_47656_125 = 1'h1;
  assign T_47656_126 = 1'h1;
  assign T_47656_127 = 1'h1;
  assign T_47656_128 = 1'h1;
  assign T_47656_129 = 1'h1;
  assign T_47656_130 = 1'h1;
  assign T_47656_131 = 1'h1;
  assign T_47656_132 = 1'h1;
  assign T_47656_133 = 1'h1;
  assign T_47656_134 = 1'h1;
  assign T_47656_135 = 1'h1;
  assign T_47656_136 = 1'h1;
  assign T_47656_137 = 1'h1;
  assign T_47656_138 = 1'h1;
  assign T_47656_139 = 1'h1;
  assign T_47656_140 = 1'h1;
  assign T_47656_141 = 1'h1;
  assign T_47656_142 = 1'h1;
  assign T_47656_143 = 1'h1;
  assign T_47656_144 = 1'h1;
  assign T_47656_145 = 1'h1;
  assign T_47656_146 = 1'h1;
  assign T_47656_147 = 1'h1;
  assign T_47656_148 = 1'h1;
  assign T_47656_149 = 1'h1;
  assign T_47656_150 = 1'h1;
  assign T_47656_151 = 1'h1;
  assign T_47656_152 = 1'h1;
  assign T_47656_153 = 1'h1;
  assign T_47656_154 = 1'h1;
  assign T_47656_155 = 1'h1;
  assign T_47656_156 = 1'h1;
  assign T_47656_157 = 1'h1;
  assign T_47656_158 = 1'h1;
  assign T_47656_159 = 1'h1;
  assign T_47656_160 = 1'h1;
  assign T_47656_161 = 1'h1;
  assign T_47656_162 = 1'h1;
  assign T_47656_163 = 1'h1;
  assign T_47656_164 = 1'h1;
  assign T_47656_165 = 1'h1;
  assign T_47656_166 = 1'h1;
  assign T_47656_167 = 1'h1;
  assign T_47656_168 = 1'h1;
  assign T_47656_169 = 1'h1;
  assign T_47656_170 = 1'h1;
  assign T_47656_171 = 1'h1;
  assign T_47656_172 = 1'h1;
  assign T_47656_173 = 1'h1;
  assign T_47656_174 = 1'h1;
  assign T_47656_175 = 1'h1;
  assign T_47656_176 = 1'h1;
  assign T_47656_177 = 1'h1;
  assign T_47656_178 = 1'h1;
  assign T_47656_179 = 1'h1;
  assign T_47656_180 = 1'h1;
  assign T_47656_181 = 1'h1;
  assign T_47656_182 = 1'h1;
  assign T_47656_183 = 1'h1;
  assign T_47656_184 = 1'h1;
  assign T_47656_185 = 1'h1;
  assign T_47656_186 = 1'h1;
  assign T_47656_187 = 1'h1;
  assign T_47656_188 = 1'h1;
  assign T_47656_189 = 1'h1;
  assign T_47656_190 = 1'h1;
  assign T_47656_191 = 1'h1;
  assign T_47656_192 = 1'h1;
  assign T_47656_193 = 1'h1;
  assign T_47656_194 = 1'h1;
  assign T_47656_195 = 1'h1;
  assign T_47656_196 = 1'h1;
  assign T_47656_197 = 1'h1;
  assign T_47656_198 = 1'h1;
  assign T_47656_199 = 1'h1;
  assign T_47656_200 = 1'h1;
  assign T_47656_201 = 1'h1;
  assign T_47656_202 = 1'h1;
  assign T_47656_203 = 1'h1;
  assign T_47656_204 = 1'h1;
  assign T_47656_205 = 1'h1;
  assign T_47656_206 = 1'h1;
  assign T_47656_207 = 1'h1;
  assign T_47656_208 = 1'h1;
  assign T_47656_209 = 1'h1;
  assign T_47656_210 = 1'h1;
  assign T_47656_211 = 1'h1;
  assign T_47656_212 = 1'h1;
  assign T_47656_213 = 1'h1;
  assign T_47656_214 = 1'h1;
  assign T_47656_215 = 1'h1;
  assign T_47656_216 = 1'h1;
  assign T_47656_217 = 1'h1;
  assign T_47656_218 = 1'h1;
  assign T_47656_219 = 1'h1;
  assign T_47656_220 = 1'h1;
  assign T_47656_221 = 1'h1;
  assign T_47656_222 = 1'h1;
  assign T_47656_223 = 1'h1;
  assign T_47656_224 = 1'h1;
  assign T_47656_225 = 1'h1;
  assign T_47656_226 = 1'h1;
  assign T_47656_227 = 1'h1;
  assign T_47656_228 = 1'h1;
  assign T_47656_229 = 1'h1;
  assign T_47656_230 = 1'h1;
  assign T_47656_231 = 1'h1;
  assign T_47656_232 = 1'h1;
  assign T_47656_233 = 1'h1;
  assign T_47656_234 = 1'h1;
  assign T_47656_235 = 1'h1;
  assign T_47656_236 = 1'h1;
  assign T_47656_237 = 1'h1;
  assign T_47656_238 = 1'h1;
  assign T_47656_239 = 1'h1;
  assign T_47656_240 = 1'h1;
  assign T_47656_241 = 1'h1;
  assign T_47656_242 = 1'h1;
  assign T_47656_243 = 1'h1;
  assign T_47656_244 = 1'h1;
  assign T_47656_245 = 1'h1;
  assign T_47656_246 = 1'h1;
  assign T_47656_247 = 1'h1;
  assign T_47656_248 = 1'h1;
  assign T_47656_249 = 1'h1;
  assign T_47656_250 = 1'h1;
  assign T_47656_251 = 1'h1;
  assign T_47656_252 = 1'h1;
  assign T_47656_253 = 1'h1;
  assign T_47656_254 = 1'h1;
  assign T_47656_255 = 1'h1;
  assign T_47656_256 = 1'h1;
  assign T_47656_257 = 1'h1;
  assign T_47656_258 = 1'h1;
  assign T_47656_259 = 1'h1;
  assign T_47656_260 = 1'h1;
  assign T_47656_261 = 1'h1;
  assign T_47656_262 = 1'h1;
  assign T_47656_263 = 1'h1;
  assign T_47656_264 = 1'h1;
  assign T_47656_265 = 1'h1;
  assign T_47656_266 = 1'h1;
  assign T_47656_267 = 1'h1;
  assign T_47656_268 = 1'h1;
  assign T_47656_269 = 1'h1;
  assign T_47656_270 = 1'h1;
  assign T_47656_271 = 1'h1;
  assign T_47656_272 = 1'h1;
  assign T_47656_273 = 1'h1;
  assign T_47656_274 = 1'h1;
  assign T_47656_275 = 1'h1;
  assign T_47656_276 = 1'h1;
  assign T_47656_277 = 1'h1;
  assign T_47656_278 = 1'h1;
  assign T_47656_279 = 1'h1;
  assign T_47656_280 = 1'h1;
  assign T_47656_281 = 1'h1;
  assign T_47656_282 = 1'h1;
  assign T_47656_283 = 1'h1;
  assign T_47656_284 = 1'h1;
  assign T_47656_285 = 1'h1;
  assign T_47656_286 = 1'h1;
  assign T_47656_287 = 1'h1;
  assign T_47656_288 = 1'h1;
  assign T_47656_289 = 1'h1;
  assign T_47656_290 = 1'h1;
  assign T_47656_291 = 1'h1;
  assign T_47656_292 = 1'h1;
  assign T_47656_293 = 1'h1;
  assign T_47656_294 = 1'h1;
  assign T_47656_295 = 1'h1;
  assign T_47656_296 = 1'h1;
  assign T_47656_297 = 1'h1;
  assign T_47656_298 = 1'h1;
  assign T_47656_299 = 1'h1;
  assign T_47656_300 = 1'h1;
  assign T_47656_301 = 1'h1;
  assign T_47656_302 = 1'h1;
  assign T_47656_303 = 1'h1;
  assign T_47656_304 = 1'h1;
  assign T_47656_305 = 1'h1;
  assign T_47656_306 = 1'h1;
  assign T_47656_307 = 1'h1;
  assign T_47656_308 = 1'h1;
  assign T_47656_309 = 1'h1;
  assign T_47656_310 = 1'h1;
  assign T_47656_311 = 1'h1;
  assign T_47656_312 = 1'h1;
  assign T_47656_313 = 1'h1;
  assign T_47656_314 = 1'h1;
  assign T_47656_315 = 1'h1;
  assign T_47656_316 = 1'h1;
  assign T_47656_317 = 1'h1;
  assign T_47656_318 = 1'h1;
  assign T_47656_319 = 1'h1;
  assign T_47656_320 = 1'h1;
  assign T_47656_321 = 1'h1;
  assign T_47656_322 = 1'h1;
  assign T_47656_323 = 1'h1;
  assign T_47656_324 = 1'h1;
  assign T_47656_325 = 1'h1;
  assign T_47656_326 = 1'h1;
  assign T_47656_327 = 1'h1;
  assign T_47656_328 = 1'h1;
  assign T_47656_329 = 1'h1;
  assign T_47656_330 = 1'h1;
  assign T_47656_331 = 1'h1;
  assign T_47656_332 = 1'h1;
  assign T_47656_333 = 1'h1;
  assign T_47656_334 = 1'h1;
  assign T_47656_335 = 1'h1;
  assign T_47656_336 = 1'h1;
  assign T_47656_337 = 1'h1;
  assign T_47656_338 = 1'h1;
  assign T_47656_339 = 1'h1;
  assign T_47656_340 = 1'h1;
  assign T_47656_341 = 1'h1;
  assign T_47656_342 = 1'h1;
  assign T_47656_343 = 1'h1;
  assign T_47656_344 = 1'h1;
  assign T_47656_345 = 1'h1;
  assign T_47656_346 = 1'h1;
  assign T_47656_347 = 1'h1;
  assign T_47656_348 = 1'h1;
  assign T_47656_349 = 1'h1;
  assign T_47656_350 = 1'h1;
  assign T_47656_351 = 1'h1;
  assign T_47656_352 = 1'h1;
  assign T_47656_353 = 1'h1;
  assign T_47656_354 = 1'h1;
  assign T_47656_355 = 1'h1;
  assign T_47656_356 = 1'h1;
  assign T_47656_357 = 1'h1;
  assign T_47656_358 = 1'h1;
  assign T_47656_359 = 1'h1;
  assign T_47656_360 = 1'h1;
  assign T_47656_361 = 1'h1;
  assign T_47656_362 = 1'h1;
  assign T_47656_363 = 1'h1;
  assign T_47656_364 = 1'h1;
  assign T_47656_365 = 1'h1;
  assign T_47656_366 = 1'h1;
  assign T_47656_367 = 1'h1;
  assign T_47656_368 = 1'h1;
  assign T_47656_369 = 1'h1;
  assign T_47656_370 = 1'h1;
  assign T_47656_371 = 1'h1;
  assign T_47656_372 = 1'h1;
  assign T_47656_373 = 1'h1;
  assign T_47656_374 = 1'h1;
  assign T_47656_375 = 1'h1;
  assign T_47656_376 = 1'h1;
  assign T_47656_377 = 1'h1;
  assign T_47656_378 = 1'h1;
  assign T_47656_379 = 1'h1;
  assign T_47656_380 = 1'h1;
  assign T_47656_381 = 1'h1;
  assign T_47656_382 = 1'h1;
  assign T_47656_383 = 1'h1;
  assign T_47656_384 = 1'h1;
  assign T_47656_385 = 1'h1;
  assign T_47656_386 = 1'h1;
  assign T_47656_387 = 1'h1;
  assign T_47656_388 = 1'h1;
  assign T_47656_389 = 1'h1;
  assign T_47656_390 = 1'h1;
  assign T_47656_391 = 1'h1;
  assign T_47656_392 = 1'h1;
  assign T_47656_393 = 1'h1;
  assign T_47656_394 = 1'h1;
  assign T_47656_395 = 1'h1;
  assign T_47656_396 = 1'h1;
  assign T_47656_397 = 1'h1;
  assign T_47656_398 = 1'h1;
  assign T_47656_399 = 1'h1;
  assign T_47656_400 = 1'h1;
  assign T_47656_401 = 1'h1;
  assign T_47656_402 = 1'h1;
  assign T_47656_403 = 1'h1;
  assign T_47656_404 = 1'h1;
  assign T_47656_405 = 1'h1;
  assign T_47656_406 = 1'h1;
  assign T_47656_407 = 1'h1;
  assign T_47656_408 = 1'h1;
  assign T_47656_409 = 1'h1;
  assign T_47656_410 = 1'h1;
  assign T_47656_411 = 1'h1;
  assign T_47656_412 = 1'h1;
  assign T_47656_413 = 1'h1;
  assign T_47656_414 = 1'h1;
  assign T_47656_415 = 1'h1;
  assign T_47656_416 = 1'h1;
  assign T_47656_417 = 1'h1;
  assign T_47656_418 = 1'h1;
  assign T_47656_419 = 1'h1;
  assign T_47656_420 = 1'h1;
  assign T_47656_421 = 1'h1;
  assign T_47656_422 = 1'h1;
  assign T_47656_423 = 1'h1;
  assign T_47656_424 = 1'h1;
  assign T_47656_425 = 1'h1;
  assign T_47656_426 = 1'h1;
  assign T_47656_427 = 1'h1;
  assign T_47656_428 = 1'h1;
  assign T_47656_429 = 1'h1;
  assign T_47656_430 = 1'h1;
  assign T_47656_431 = 1'h1;
  assign T_47656_432 = 1'h1;
  assign T_47656_433 = 1'h1;
  assign T_47656_434 = 1'h1;
  assign T_47656_435 = 1'h1;
  assign T_47656_436 = 1'h1;
  assign T_47656_437 = 1'h1;
  assign T_47656_438 = 1'h1;
  assign T_47656_439 = 1'h1;
  assign T_47656_440 = 1'h1;
  assign T_47656_441 = 1'h1;
  assign T_47656_442 = 1'h1;
  assign T_47656_443 = 1'h1;
  assign T_47656_444 = 1'h1;
  assign T_47656_445 = 1'h1;
  assign T_47656_446 = 1'h1;
  assign T_47656_447 = 1'h1;
  assign T_47656_448 = 1'h1;
  assign T_47656_449 = 1'h1;
  assign T_47656_450 = 1'h1;
  assign T_47656_451 = 1'h1;
  assign T_47656_452 = 1'h1;
  assign T_47656_453 = 1'h1;
  assign T_47656_454 = 1'h1;
  assign T_47656_455 = 1'h1;
  assign T_47656_456 = 1'h1;
  assign T_47656_457 = 1'h1;
  assign T_47656_458 = 1'h1;
  assign T_47656_459 = 1'h1;
  assign T_47656_460 = 1'h1;
  assign T_47656_461 = 1'h1;
  assign T_47656_462 = 1'h1;
  assign T_47656_463 = 1'h1;
  assign T_47656_464 = 1'h1;
  assign T_47656_465 = 1'h1;
  assign T_47656_466 = 1'h1;
  assign T_47656_467 = 1'h1;
  assign T_47656_468 = 1'h1;
  assign T_47656_469 = 1'h1;
  assign T_47656_470 = 1'h1;
  assign T_47656_471 = 1'h1;
  assign T_47656_472 = 1'h1;
  assign T_47656_473 = 1'h1;
  assign T_47656_474 = 1'h1;
  assign T_47656_475 = 1'h1;
  assign T_47656_476 = 1'h1;
  assign T_47656_477 = 1'h1;
  assign T_47656_478 = 1'h1;
  assign T_47656_479 = 1'h1;
  assign T_47656_480 = 1'h1;
  assign T_47656_481 = 1'h1;
  assign T_47656_482 = 1'h1;
  assign T_47656_483 = 1'h1;
  assign T_47656_484 = 1'h1;
  assign T_47656_485 = 1'h1;
  assign T_47656_486 = 1'h1;
  assign T_47656_487 = 1'h1;
  assign T_47656_488 = 1'h1;
  assign T_47656_489 = 1'h1;
  assign T_47656_490 = 1'h1;
  assign T_47656_491 = 1'h1;
  assign T_47656_492 = 1'h1;
  assign T_47656_493 = 1'h1;
  assign T_47656_494 = 1'h1;
  assign T_47656_495 = 1'h1;
  assign T_47656_496 = 1'h1;
  assign T_47656_497 = 1'h1;
  assign T_47656_498 = 1'h1;
  assign T_47656_499 = 1'h1;
  assign T_47656_500 = 1'h1;
  assign T_47656_501 = 1'h1;
  assign T_47656_502 = 1'h1;
  assign T_47656_503 = 1'h1;
  assign T_47656_504 = 1'h1;
  assign T_47656_505 = 1'h1;
  assign T_47656_506 = 1'h1;
  assign T_47656_507 = 1'h1;
  assign T_47656_508 = 1'h1;
  assign T_47656_509 = 1'h1;
  assign T_47656_510 = 1'h1;
  assign T_47656_511 = 1'h1;
  assign T_48687_0 = T_8270;
  assign T_48687_1 = T_9573;
  assign T_48687_2 = T_9933;
  assign T_48687_3 = T_11733;
  assign T_48687_4 = T_13213;
  assign T_48687_5 = T_8310;
  assign T_48687_6 = T_9613;
  assign T_48687_7 = T_11653;
  assign T_48687_8 = T_13013;
  assign T_48687_9 = T_9813;
  assign T_48687_10 = T_8350;
  assign T_48687_11 = T_12813;
  assign T_48687_12 = T_11573;
  assign T_48687_13 = T_9853;
  assign T_48687_14 = T_8550;
  assign T_48687_15 = T_13293;
  assign T_48687_16 = T_12733;
  assign T_48687_17 = T_10093;
  assign T_48687_18 = T_12653;
  assign T_48687_19 = T_13173;
  assign T_48687_20 = T_8590;
  assign T_48687_21 = T_9733;
  assign T_48687_22 = T_11453;
  assign T_48687_23 = T_12973;
  assign T_48687_24 = T_8430;
  assign T_48687_25 = T_8510;
  assign T_48687_26 = T_12933;
  assign T_48687_27 = T_11533;
  assign T_48687_28 = T_9653;
  assign T_48687_29 = T_9470;
  assign T_48687_30 = T_13093;
  assign T_48687_31 = T_12773;
  assign T_48687_32 = T_9973;
  assign T_48687_33 = T_9773;
  assign T_48687_34 = T_10013;
  assign T_48687_35 = T_11773;
  assign T_48687_36 = T_13053;
  assign T_48687_37 = T_8470;
  assign T_48687_38 = T_9693;
  assign T_48687_39 = T_11693;
  assign T_48687_40 = T_12893;
  assign T_48687_41 = T_9893;
  assign T_48687_42 = T_8390;
  assign T_48687_43 = T_12853;
  assign T_48687_44 = T_11493;
  assign T_48687_45 = T_10053;
  assign T_48687_46 = T_9430;
  assign T_48687_47 = T_13253;
  assign T_48687_48 = T_11813;
  assign T_48687_49 = T_11613;
  assign T_48687_50 = T_12693;
  assign T_48687_51 = T_13133;
  assign T_48687_52 = 32'h0;
  assign T_48687_53 = 32'h0;
  assign T_48687_54 = 32'h0;
  assign T_48687_55 = 32'h0;
  assign T_48687_56 = 32'h0;
  assign T_48687_57 = 32'h0;
  assign T_48687_58 = 32'h0;
  assign T_48687_59 = 32'h0;
  assign T_48687_60 = 32'h0;
  assign T_48687_61 = 32'h0;
  assign T_48687_62 = 32'h0;
  assign T_48687_63 = 32'h0;
  assign T_48687_64 = T_8231;
  assign T_48687_65 = {{12'd0}, T_12614};
  assign T_48687_66 = 32'h0;
  assign T_48687_67 = 32'h0;
  assign T_48687_68 = 32'h0;
  assign T_48687_69 = 32'h0;
  assign T_48687_70 = 32'h0;
  assign T_48687_71 = 32'h0;
  assign T_48687_72 = 32'h0;
  assign T_48687_73 = 32'h0;
  assign T_48687_74 = 32'h0;
  assign T_48687_75 = 32'h0;
  assign T_48687_76 = 32'h0;
  assign T_48687_77 = 32'h0;
  assign T_48687_78 = 32'h0;
  assign T_48687_79 = 32'h0;
  assign T_48687_80 = 32'h0;
  assign T_48687_81 = 32'h0;
  assign T_48687_82 = 32'h0;
  assign T_48687_83 = 32'h0;
  assign T_48687_84 = 32'h0;
  assign T_48687_85 = 32'h0;
  assign T_48687_86 = 32'h0;
  assign T_48687_87 = 32'h0;
  assign T_48687_88 = 32'h0;
  assign T_48687_89 = 32'h0;
  assign T_48687_90 = 32'h0;
  assign T_48687_91 = 32'h0;
  assign T_48687_92 = 32'h0;
  assign T_48687_93 = 32'h0;
  assign T_48687_94 = 32'h0;
  assign T_48687_95 = 32'h0;
  assign T_48687_96 = 32'h0;
  assign T_48687_97 = 32'h0;
  assign T_48687_98 = 32'h0;
  assign T_48687_99 = 32'h0;
  assign T_48687_100 = 32'h0;
  assign T_48687_101 = 32'h0;
  assign T_48687_102 = 32'h0;
  assign T_48687_103 = 32'h0;
  assign T_48687_104 = 32'h0;
  assign T_48687_105 = 32'h0;
  assign T_48687_106 = 32'h0;
  assign T_48687_107 = 32'h0;
  assign T_48687_108 = 32'h0;
  assign T_48687_109 = 32'h0;
  assign T_48687_110 = 32'h0;
  assign T_48687_111 = 32'h0;
  assign T_48687_112 = 32'h0;
  assign T_48687_113 = 32'h0;
  assign T_48687_114 = 32'h0;
  assign T_48687_115 = 32'h0;
  assign T_48687_116 = 32'h0;
  assign T_48687_117 = 32'h0;
  assign T_48687_118 = 32'h0;
  assign T_48687_119 = 32'h0;
  assign T_48687_120 = 32'h0;
  assign T_48687_121 = 32'h0;
  assign T_48687_122 = 32'h0;
  assign T_48687_123 = 32'h0;
  assign T_48687_124 = 32'h0;
  assign T_48687_125 = 32'h0;
  assign T_48687_126 = 32'h0;
  assign T_48687_127 = 32'h0;
  assign T_48687_128 = T_11414;
  assign T_48687_129 = {{12'd0}, T_9391};
  assign T_48687_130 = 32'h0;
  assign T_48687_131 = 32'h0;
  assign T_48687_132 = 32'h0;
  assign T_48687_133 = 32'h0;
  assign T_48687_134 = 32'h0;
  assign T_48687_135 = 32'h0;
  assign T_48687_136 = 32'h0;
  assign T_48687_137 = 32'h0;
  assign T_48687_138 = 32'h0;
  assign T_48687_139 = 32'h0;
  assign T_48687_140 = 32'h0;
  assign T_48687_141 = 32'h0;
  assign T_48687_142 = 32'h0;
  assign T_48687_143 = 32'h0;
  assign T_48687_144 = 32'h0;
  assign T_48687_145 = 32'h0;
  assign T_48687_146 = 32'h0;
  assign T_48687_147 = 32'h0;
  assign T_48687_148 = 32'h0;
  assign T_48687_149 = 32'h0;
  assign T_48687_150 = 32'h0;
  assign T_48687_151 = 32'h0;
  assign T_48687_152 = 32'h0;
  assign T_48687_153 = 32'h0;
  assign T_48687_154 = 32'h0;
  assign T_48687_155 = 32'h0;
  assign T_48687_156 = 32'h0;
  assign T_48687_157 = 32'h0;
  assign T_48687_158 = 32'h0;
  assign T_48687_159 = 32'h0;
  assign T_48687_160 = 32'h0;
  assign T_48687_161 = 32'h0;
  assign T_48687_162 = 32'h0;
  assign T_48687_163 = 32'h0;
  assign T_48687_164 = 32'h0;
  assign T_48687_165 = 32'h0;
  assign T_48687_166 = 32'h0;
  assign T_48687_167 = 32'h0;
  assign T_48687_168 = 32'h0;
  assign T_48687_169 = 32'h0;
  assign T_48687_170 = 32'h0;
  assign T_48687_171 = 32'h0;
  assign T_48687_172 = 32'h0;
  assign T_48687_173 = 32'h0;
  assign T_48687_174 = 32'h0;
  assign T_48687_175 = 32'h0;
  assign T_48687_176 = 32'h0;
  assign T_48687_177 = 32'h0;
  assign T_48687_178 = 32'h0;
  assign T_48687_179 = 32'h0;
  assign T_48687_180 = 32'h0;
  assign T_48687_181 = 32'h0;
  assign T_48687_182 = 32'h0;
  assign T_48687_183 = 32'h0;
  assign T_48687_184 = 32'h0;
  assign T_48687_185 = 32'h0;
  assign T_48687_186 = 32'h0;
  assign T_48687_187 = 32'h0;
  assign T_48687_188 = 32'h0;
  assign T_48687_189 = 32'h0;
  assign T_48687_190 = 32'h0;
  assign T_48687_191 = 32'h0;
  assign T_48687_192 = 32'h0;
  assign T_48687_193 = 32'h0;
  assign T_48687_194 = 32'h0;
  assign T_48687_195 = 32'h0;
  assign T_48687_196 = 32'h0;
  assign T_48687_197 = 32'h0;
  assign T_48687_198 = 32'h0;
  assign T_48687_199 = 32'h0;
  assign T_48687_200 = 32'h0;
  assign T_48687_201 = 32'h0;
  assign T_48687_202 = 32'h0;
  assign T_48687_203 = 32'h0;
  assign T_48687_204 = 32'h0;
  assign T_48687_205 = 32'h0;
  assign T_48687_206 = 32'h0;
  assign T_48687_207 = 32'h0;
  assign T_48687_208 = 32'h0;
  assign T_48687_209 = 32'h0;
  assign T_48687_210 = 32'h0;
  assign T_48687_211 = 32'h0;
  assign T_48687_212 = 32'h0;
  assign T_48687_213 = 32'h0;
  assign T_48687_214 = 32'h0;
  assign T_48687_215 = 32'h0;
  assign T_48687_216 = 32'h0;
  assign T_48687_217 = 32'h0;
  assign T_48687_218 = 32'h0;
  assign T_48687_219 = 32'h0;
  assign T_48687_220 = 32'h0;
  assign T_48687_221 = 32'h0;
  assign T_48687_222 = 32'h0;
  assign T_48687_223 = 32'h0;
  assign T_48687_224 = 32'h0;
  assign T_48687_225 = 32'h0;
  assign T_48687_226 = 32'h0;
  assign T_48687_227 = 32'h0;
  assign T_48687_228 = 32'h0;
  assign T_48687_229 = 32'h0;
  assign T_48687_230 = 32'h0;
  assign T_48687_231 = 32'h0;
  assign T_48687_232 = 32'h0;
  assign T_48687_233 = 32'h0;
  assign T_48687_234 = 32'h0;
  assign T_48687_235 = 32'h0;
  assign T_48687_236 = 32'h0;
  assign T_48687_237 = 32'h0;
  assign T_48687_238 = 32'h0;
  assign T_48687_239 = 32'h0;
  assign T_48687_240 = 32'h0;
  assign T_48687_241 = 32'h0;
  assign T_48687_242 = 32'h0;
  assign T_48687_243 = 32'h0;
  assign T_48687_244 = 32'h0;
  assign T_48687_245 = 32'h0;
  assign T_48687_246 = 32'h0;
  assign T_48687_247 = 32'h0;
  assign T_48687_248 = 32'h0;
  assign T_48687_249 = 32'h0;
  assign T_48687_250 = 32'h0;
  assign T_48687_251 = 32'h0;
  assign T_48687_252 = 32'h0;
  assign T_48687_253 = 32'h0;
  assign T_48687_254 = 32'h0;
  assign T_48687_255 = 32'h0;
  assign T_48687_256 = T_10133;
  assign T_48687_257 = T_9533;
  assign T_48687_258 = 32'h0;
  assign T_48687_259 = 32'h0;
  assign T_48687_260 = 32'h0;
  assign T_48687_261 = 32'h0;
  assign T_48687_262 = 32'h0;
  assign T_48687_263 = 32'h0;
  assign T_48687_264 = 32'h0;
  assign T_48687_265 = 32'h0;
  assign T_48687_266 = 32'h0;
  assign T_48687_267 = 32'h0;
  assign T_48687_268 = 32'h0;
  assign T_48687_269 = 32'h0;
  assign T_48687_270 = 32'h0;
  assign T_48687_271 = 32'h0;
  assign T_48687_272 = 32'h0;
  assign T_48687_273 = 32'h0;
  assign T_48687_274 = 32'h0;
  assign T_48687_275 = 32'h0;
  assign T_48687_276 = 32'h0;
  assign T_48687_277 = 32'h0;
  assign T_48687_278 = 32'h0;
  assign T_48687_279 = 32'h0;
  assign T_48687_280 = 32'h0;
  assign T_48687_281 = 32'h0;
  assign T_48687_282 = 32'h0;
  assign T_48687_283 = 32'h0;
  assign T_48687_284 = 32'h0;
  assign T_48687_285 = 32'h0;
  assign T_48687_286 = 32'h0;
  assign T_48687_287 = 32'h0;
  assign T_48687_288 = 32'h0;
  assign T_48687_289 = 32'h0;
  assign T_48687_290 = 32'h0;
  assign T_48687_291 = 32'h0;
  assign T_48687_292 = 32'h0;
  assign T_48687_293 = 32'h0;
  assign T_48687_294 = 32'h0;
  assign T_48687_295 = 32'h0;
  assign T_48687_296 = 32'h0;
  assign T_48687_297 = 32'h0;
  assign T_48687_298 = 32'h0;
  assign T_48687_299 = 32'h0;
  assign T_48687_300 = 32'h0;
  assign T_48687_301 = 32'h0;
  assign T_48687_302 = 32'h0;
  assign T_48687_303 = 32'h0;
  assign T_48687_304 = 32'h0;
  assign T_48687_305 = 32'h0;
  assign T_48687_306 = 32'h0;
  assign T_48687_307 = 32'h0;
  assign T_48687_308 = 32'h0;
  assign T_48687_309 = 32'h0;
  assign T_48687_310 = 32'h0;
  assign T_48687_311 = 32'h0;
  assign T_48687_312 = 32'h0;
  assign T_48687_313 = 32'h0;
  assign T_48687_314 = 32'h0;
  assign T_48687_315 = 32'h0;
  assign T_48687_316 = 32'h0;
  assign T_48687_317 = 32'h0;
  assign T_48687_318 = 32'h0;
  assign T_48687_319 = 32'h0;
  assign T_48687_320 = 32'h0;
  assign T_48687_321 = 32'h0;
  assign T_48687_322 = 32'h0;
  assign T_48687_323 = 32'h0;
  assign T_48687_324 = 32'h0;
  assign T_48687_325 = 32'h0;
  assign T_48687_326 = 32'h0;
  assign T_48687_327 = 32'h0;
  assign T_48687_328 = 32'h0;
  assign T_48687_329 = 32'h0;
  assign T_48687_330 = 32'h0;
  assign T_48687_331 = 32'h0;
  assign T_48687_332 = 32'h0;
  assign T_48687_333 = 32'h0;
  assign T_48687_334 = 32'h0;
  assign T_48687_335 = 32'h0;
  assign T_48687_336 = 32'h0;
  assign T_48687_337 = 32'h0;
  assign T_48687_338 = 32'h0;
  assign T_48687_339 = 32'h0;
  assign T_48687_340 = 32'h0;
  assign T_48687_341 = 32'h0;
  assign T_48687_342 = 32'h0;
  assign T_48687_343 = 32'h0;
  assign T_48687_344 = 32'h0;
  assign T_48687_345 = 32'h0;
  assign T_48687_346 = 32'h0;
  assign T_48687_347 = 32'h0;
  assign T_48687_348 = 32'h0;
  assign T_48687_349 = 32'h0;
  assign T_48687_350 = 32'h0;
  assign T_48687_351 = 32'h0;
  assign T_48687_352 = 32'h0;
  assign T_48687_353 = 32'h0;
  assign T_48687_354 = 32'h0;
  assign T_48687_355 = 32'h0;
  assign T_48687_356 = 32'h0;
  assign T_48687_357 = 32'h0;
  assign T_48687_358 = 32'h0;
  assign T_48687_359 = 32'h0;
  assign T_48687_360 = 32'h0;
  assign T_48687_361 = 32'h0;
  assign T_48687_362 = 32'h0;
  assign T_48687_363 = 32'h0;
  assign T_48687_364 = 32'h0;
  assign T_48687_365 = 32'h0;
  assign T_48687_366 = 32'h0;
  assign T_48687_367 = 32'h0;
  assign T_48687_368 = 32'h0;
  assign T_48687_369 = 32'h0;
  assign T_48687_370 = 32'h0;
  assign T_48687_371 = 32'h0;
  assign T_48687_372 = 32'h0;
  assign T_48687_373 = 32'h0;
  assign T_48687_374 = 32'h0;
  assign T_48687_375 = 32'h0;
  assign T_48687_376 = 32'h0;
  assign T_48687_377 = 32'h0;
  assign T_48687_378 = 32'h0;
  assign T_48687_379 = 32'h0;
  assign T_48687_380 = 32'h0;
  assign T_48687_381 = 32'h0;
  assign T_48687_382 = 32'h0;
  assign T_48687_383 = 32'h0;
  assign T_48687_384 = 32'h0;
  assign T_48687_385 = 32'h0;
  assign T_48687_386 = 32'h0;
  assign T_48687_387 = 32'h0;
  assign T_48687_388 = 32'h0;
  assign T_48687_389 = 32'h0;
  assign T_48687_390 = 32'h0;
  assign T_48687_391 = 32'h0;
  assign T_48687_392 = 32'h0;
  assign T_48687_393 = 32'h0;
  assign T_48687_394 = 32'h0;
  assign T_48687_395 = 32'h0;
  assign T_48687_396 = 32'h0;
  assign T_48687_397 = 32'h0;
  assign T_48687_398 = 32'h0;
  assign T_48687_399 = 32'h0;
  assign T_48687_400 = 32'h0;
  assign T_48687_401 = 32'h0;
  assign T_48687_402 = 32'h0;
  assign T_48687_403 = 32'h0;
  assign T_48687_404 = 32'h0;
  assign T_48687_405 = 32'h0;
  assign T_48687_406 = 32'h0;
  assign T_48687_407 = 32'h0;
  assign T_48687_408 = 32'h0;
  assign T_48687_409 = 32'h0;
  assign T_48687_410 = 32'h0;
  assign T_48687_411 = 32'h0;
  assign T_48687_412 = 32'h0;
  assign T_48687_413 = 32'h0;
  assign T_48687_414 = 32'h0;
  assign T_48687_415 = 32'h0;
  assign T_48687_416 = 32'h0;
  assign T_48687_417 = 32'h0;
  assign T_48687_418 = 32'h0;
  assign T_48687_419 = 32'h0;
  assign T_48687_420 = 32'h0;
  assign T_48687_421 = 32'h0;
  assign T_48687_422 = 32'h0;
  assign T_48687_423 = 32'h0;
  assign T_48687_424 = 32'h0;
  assign T_48687_425 = 32'h0;
  assign T_48687_426 = 32'h0;
  assign T_48687_427 = 32'h0;
  assign T_48687_428 = 32'h0;
  assign T_48687_429 = 32'h0;
  assign T_48687_430 = 32'h0;
  assign T_48687_431 = 32'h0;
  assign T_48687_432 = 32'h0;
  assign T_48687_433 = 32'h0;
  assign T_48687_434 = 32'h0;
  assign T_48687_435 = 32'h0;
  assign T_48687_436 = 32'h0;
  assign T_48687_437 = 32'h0;
  assign T_48687_438 = 32'h0;
  assign T_48687_439 = 32'h0;
  assign T_48687_440 = 32'h0;
  assign T_48687_441 = 32'h0;
  assign T_48687_442 = 32'h0;
  assign T_48687_443 = 32'h0;
  assign T_48687_444 = 32'h0;
  assign T_48687_445 = 32'h0;
  assign T_48687_446 = 32'h0;
  assign T_48687_447 = 32'h0;
  assign T_48687_448 = 32'h0;
  assign T_48687_449 = 32'h0;
  assign T_48687_450 = 32'h0;
  assign T_48687_451 = 32'h0;
  assign T_48687_452 = 32'h0;
  assign T_48687_453 = 32'h0;
  assign T_48687_454 = 32'h0;
  assign T_48687_455 = 32'h0;
  assign T_48687_456 = 32'h0;
  assign T_48687_457 = 32'h0;
  assign T_48687_458 = 32'h0;
  assign T_48687_459 = 32'h0;
  assign T_48687_460 = 32'h0;
  assign T_48687_461 = 32'h0;
  assign T_48687_462 = 32'h0;
  assign T_48687_463 = 32'h0;
  assign T_48687_464 = 32'h0;
  assign T_48687_465 = 32'h0;
  assign T_48687_466 = 32'h0;
  assign T_48687_467 = 32'h0;
  assign T_48687_468 = 32'h0;
  assign T_48687_469 = 32'h0;
  assign T_48687_470 = 32'h0;
  assign T_48687_471 = 32'h0;
  assign T_48687_472 = 32'h0;
  assign T_48687_473 = 32'h0;
  assign T_48687_474 = 32'h0;
  assign T_48687_475 = 32'h0;
  assign T_48687_476 = 32'h0;
  assign T_48687_477 = 32'h0;
  assign T_48687_478 = 32'h0;
  assign T_48687_479 = 32'h0;
  assign T_48687_480 = 32'h0;
  assign T_48687_481 = 32'h0;
  assign T_48687_482 = 32'h0;
  assign T_48687_483 = 32'h0;
  assign T_48687_484 = 32'h0;
  assign T_48687_485 = 32'h0;
  assign T_48687_486 = 32'h0;
  assign T_48687_487 = 32'h0;
  assign T_48687_488 = 32'h0;
  assign T_48687_489 = 32'h0;
  assign T_48687_490 = 32'h0;
  assign T_48687_491 = 32'h0;
  assign T_48687_492 = 32'h0;
  assign T_48687_493 = 32'h0;
  assign T_48687_494 = 32'h0;
  assign T_48687_495 = 32'h0;
  assign T_48687_496 = 32'h0;
  assign T_48687_497 = 32'h0;
  assign T_48687_498 = 32'h0;
  assign T_48687_499 = 32'h0;
  assign T_48687_500 = 32'h0;
  assign T_48687_501 = 32'h0;
  assign T_48687_502 = 32'h0;
  assign T_48687_503 = 32'h0;
  assign T_48687_504 = 32'h0;
  assign T_48687_505 = 32'h0;
  assign T_48687_506 = 32'h0;
  assign T_48687_507 = 32'h0;
  assign T_48687_508 = 32'h0;
  assign T_48687_509 = 32'h0;
  assign T_48687_510 = 32'h0;
  assign T_48687_511 = 32'h0;
  assign GEN_7 = GEN_2977;
  assign GEN_2467 = 9'h1 == T_24222 ? T_47656_1 : T_47656_0;
  assign GEN_2468 = 9'h2 == T_24222 ? T_47656_2 : GEN_2467;
  assign GEN_2469 = 9'h3 == T_24222 ? T_47656_3 : GEN_2468;
  assign GEN_2470 = 9'h4 == T_24222 ? T_47656_4 : GEN_2469;
  assign GEN_2471 = 9'h5 == T_24222 ? T_47656_5 : GEN_2470;
  assign GEN_2472 = 9'h6 == T_24222 ? T_47656_6 : GEN_2471;
  assign GEN_2473 = 9'h7 == T_24222 ? T_47656_7 : GEN_2472;
  assign GEN_2474 = 9'h8 == T_24222 ? T_47656_8 : GEN_2473;
  assign GEN_2475 = 9'h9 == T_24222 ? T_47656_9 : GEN_2474;
  assign GEN_2476 = 9'ha == T_24222 ? T_47656_10 : GEN_2475;
  assign GEN_2477 = 9'hb == T_24222 ? T_47656_11 : GEN_2476;
  assign GEN_2478 = 9'hc == T_24222 ? T_47656_12 : GEN_2477;
  assign GEN_2479 = 9'hd == T_24222 ? T_47656_13 : GEN_2478;
  assign GEN_2480 = 9'he == T_24222 ? T_47656_14 : GEN_2479;
  assign GEN_2481 = 9'hf == T_24222 ? T_47656_15 : GEN_2480;
  assign GEN_2482 = 9'h10 == T_24222 ? T_47656_16 : GEN_2481;
  assign GEN_2483 = 9'h11 == T_24222 ? T_47656_17 : GEN_2482;
  assign GEN_2484 = 9'h12 == T_24222 ? T_47656_18 : GEN_2483;
  assign GEN_2485 = 9'h13 == T_24222 ? T_47656_19 : GEN_2484;
  assign GEN_2486 = 9'h14 == T_24222 ? T_47656_20 : GEN_2485;
  assign GEN_2487 = 9'h15 == T_24222 ? T_47656_21 : GEN_2486;
  assign GEN_2488 = 9'h16 == T_24222 ? T_47656_22 : GEN_2487;
  assign GEN_2489 = 9'h17 == T_24222 ? T_47656_23 : GEN_2488;
  assign GEN_2490 = 9'h18 == T_24222 ? T_47656_24 : GEN_2489;
  assign GEN_2491 = 9'h19 == T_24222 ? T_47656_25 : GEN_2490;
  assign GEN_2492 = 9'h1a == T_24222 ? T_47656_26 : GEN_2491;
  assign GEN_2493 = 9'h1b == T_24222 ? T_47656_27 : GEN_2492;
  assign GEN_2494 = 9'h1c == T_24222 ? T_47656_28 : GEN_2493;
  assign GEN_2495 = 9'h1d == T_24222 ? T_47656_29 : GEN_2494;
  assign GEN_2496 = 9'h1e == T_24222 ? T_47656_30 : GEN_2495;
  assign GEN_2497 = 9'h1f == T_24222 ? T_47656_31 : GEN_2496;
  assign GEN_2498 = 9'h20 == T_24222 ? T_47656_32 : GEN_2497;
  assign GEN_2499 = 9'h21 == T_24222 ? T_47656_33 : GEN_2498;
  assign GEN_2500 = 9'h22 == T_24222 ? T_47656_34 : GEN_2499;
  assign GEN_2501 = 9'h23 == T_24222 ? T_47656_35 : GEN_2500;
  assign GEN_2502 = 9'h24 == T_24222 ? T_47656_36 : GEN_2501;
  assign GEN_2503 = 9'h25 == T_24222 ? T_47656_37 : GEN_2502;
  assign GEN_2504 = 9'h26 == T_24222 ? T_47656_38 : GEN_2503;
  assign GEN_2505 = 9'h27 == T_24222 ? T_47656_39 : GEN_2504;
  assign GEN_2506 = 9'h28 == T_24222 ? T_47656_40 : GEN_2505;
  assign GEN_2507 = 9'h29 == T_24222 ? T_47656_41 : GEN_2506;
  assign GEN_2508 = 9'h2a == T_24222 ? T_47656_42 : GEN_2507;
  assign GEN_2509 = 9'h2b == T_24222 ? T_47656_43 : GEN_2508;
  assign GEN_2510 = 9'h2c == T_24222 ? T_47656_44 : GEN_2509;
  assign GEN_2511 = 9'h2d == T_24222 ? T_47656_45 : GEN_2510;
  assign GEN_2512 = 9'h2e == T_24222 ? T_47656_46 : GEN_2511;
  assign GEN_2513 = 9'h2f == T_24222 ? T_47656_47 : GEN_2512;
  assign GEN_2514 = 9'h30 == T_24222 ? T_47656_48 : GEN_2513;
  assign GEN_2515 = 9'h31 == T_24222 ? T_47656_49 : GEN_2514;
  assign GEN_2516 = 9'h32 == T_24222 ? T_47656_50 : GEN_2515;
  assign GEN_2517 = 9'h33 == T_24222 ? T_47656_51 : GEN_2516;
  assign GEN_2518 = 9'h34 == T_24222 ? T_47656_52 : GEN_2517;
  assign GEN_2519 = 9'h35 == T_24222 ? T_47656_53 : GEN_2518;
  assign GEN_2520 = 9'h36 == T_24222 ? T_47656_54 : GEN_2519;
  assign GEN_2521 = 9'h37 == T_24222 ? T_47656_55 : GEN_2520;
  assign GEN_2522 = 9'h38 == T_24222 ? T_47656_56 : GEN_2521;
  assign GEN_2523 = 9'h39 == T_24222 ? T_47656_57 : GEN_2522;
  assign GEN_2524 = 9'h3a == T_24222 ? T_47656_58 : GEN_2523;
  assign GEN_2525 = 9'h3b == T_24222 ? T_47656_59 : GEN_2524;
  assign GEN_2526 = 9'h3c == T_24222 ? T_47656_60 : GEN_2525;
  assign GEN_2527 = 9'h3d == T_24222 ? T_47656_61 : GEN_2526;
  assign GEN_2528 = 9'h3e == T_24222 ? T_47656_62 : GEN_2527;
  assign GEN_2529 = 9'h3f == T_24222 ? T_47656_63 : GEN_2528;
  assign GEN_2530 = 9'h40 == T_24222 ? T_47656_64 : GEN_2529;
  assign GEN_2531 = 9'h41 == T_24222 ? T_47656_65 : GEN_2530;
  assign GEN_2532 = 9'h42 == T_24222 ? T_47656_66 : GEN_2531;
  assign GEN_2533 = 9'h43 == T_24222 ? T_47656_67 : GEN_2532;
  assign GEN_2534 = 9'h44 == T_24222 ? T_47656_68 : GEN_2533;
  assign GEN_2535 = 9'h45 == T_24222 ? T_47656_69 : GEN_2534;
  assign GEN_2536 = 9'h46 == T_24222 ? T_47656_70 : GEN_2535;
  assign GEN_2537 = 9'h47 == T_24222 ? T_47656_71 : GEN_2536;
  assign GEN_2538 = 9'h48 == T_24222 ? T_47656_72 : GEN_2537;
  assign GEN_2539 = 9'h49 == T_24222 ? T_47656_73 : GEN_2538;
  assign GEN_2540 = 9'h4a == T_24222 ? T_47656_74 : GEN_2539;
  assign GEN_2541 = 9'h4b == T_24222 ? T_47656_75 : GEN_2540;
  assign GEN_2542 = 9'h4c == T_24222 ? T_47656_76 : GEN_2541;
  assign GEN_2543 = 9'h4d == T_24222 ? T_47656_77 : GEN_2542;
  assign GEN_2544 = 9'h4e == T_24222 ? T_47656_78 : GEN_2543;
  assign GEN_2545 = 9'h4f == T_24222 ? T_47656_79 : GEN_2544;
  assign GEN_2546 = 9'h50 == T_24222 ? T_47656_80 : GEN_2545;
  assign GEN_2547 = 9'h51 == T_24222 ? T_47656_81 : GEN_2546;
  assign GEN_2548 = 9'h52 == T_24222 ? T_47656_82 : GEN_2547;
  assign GEN_2549 = 9'h53 == T_24222 ? T_47656_83 : GEN_2548;
  assign GEN_2550 = 9'h54 == T_24222 ? T_47656_84 : GEN_2549;
  assign GEN_2551 = 9'h55 == T_24222 ? T_47656_85 : GEN_2550;
  assign GEN_2552 = 9'h56 == T_24222 ? T_47656_86 : GEN_2551;
  assign GEN_2553 = 9'h57 == T_24222 ? T_47656_87 : GEN_2552;
  assign GEN_2554 = 9'h58 == T_24222 ? T_47656_88 : GEN_2553;
  assign GEN_2555 = 9'h59 == T_24222 ? T_47656_89 : GEN_2554;
  assign GEN_2556 = 9'h5a == T_24222 ? T_47656_90 : GEN_2555;
  assign GEN_2557 = 9'h5b == T_24222 ? T_47656_91 : GEN_2556;
  assign GEN_2558 = 9'h5c == T_24222 ? T_47656_92 : GEN_2557;
  assign GEN_2559 = 9'h5d == T_24222 ? T_47656_93 : GEN_2558;
  assign GEN_2560 = 9'h5e == T_24222 ? T_47656_94 : GEN_2559;
  assign GEN_2561 = 9'h5f == T_24222 ? T_47656_95 : GEN_2560;
  assign GEN_2562 = 9'h60 == T_24222 ? T_47656_96 : GEN_2561;
  assign GEN_2563 = 9'h61 == T_24222 ? T_47656_97 : GEN_2562;
  assign GEN_2564 = 9'h62 == T_24222 ? T_47656_98 : GEN_2563;
  assign GEN_2565 = 9'h63 == T_24222 ? T_47656_99 : GEN_2564;
  assign GEN_2566 = 9'h64 == T_24222 ? T_47656_100 : GEN_2565;
  assign GEN_2567 = 9'h65 == T_24222 ? T_47656_101 : GEN_2566;
  assign GEN_2568 = 9'h66 == T_24222 ? T_47656_102 : GEN_2567;
  assign GEN_2569 = 9'h67 == T_24222 ? T_47656_103 : GEN_2568;
  assign GEN_2570 = 9'h68 == T_24222 ? T_47656_104 : GEN_2569;
  assign GEN_2571 = 9'h69 == T_24222 ? T_47656_105 : GEN_2570;
  assign GEN_2572 = 9'h6a == T_24222 ? T_47656_106 : GEN_2571;
  assign GEN_2573 = 9'h6b == T_24222 ? T_47656_107 : GEN_2572;
  assign GEN_2574 = 9'h6c == T_24222 ? T_47656_108 : GEN_2573;
  assign GEN_2575 = 9'h6d == T_24222 ? T_47656_109 : GEN_2574;
  assign GEN_2576 = 9'h6e == T_24222 ? T_47656_110 : GEN_2575;
  assign GEN_2577 = 9'h6f == T_24222 ? T_47656_111 : GEN_2576;
  assign GEN_2578 = 9'h70 == T_24222 ? T_47656_112 : GEN_2577;
  assign GEN_2579 = 9'h71 == T_24222 ? T_47656_113 : GEN_2578;
  assign GEN_2580 = 9'h72 == T_24222 ? T_47656_114 : GEN_2579;
  assign GEN_2581 = 9'h73 == T_24222 ? T_47656_115 : GEN_2580;
  assign GEN_2582 = 9'h74 == T_24222 ? T_47656_116 : GEN_2581;
  assign GEN_2583 = 9'h75 == T_24222 ? T_47656_117 : GEN_2582;
  assign GEN_2584 = 9'h76 == T_24222 ? T_47656_118 : GEN_2583;
  assign GEN_2585 = 9'h77 == T_24222 ? T_47656_119 : GEN_2584;
  assign GEN_2586 = 9'h78 == T_24222 ? T_47656_120 : GEN_2585;
  assign GEN_2587 = 9'h79 == T_24222 ? T_47656_121 : GEN_2586;
  assign GEN_2588 = 9'h7a == T_24222 ? T_47656_122 : GEN_2587;
  assign GEN_2589 = 9'h7b == T_24222 ? T_47656_123 : GEN_2588;
  assign GEN_2590 = 9'h7c == T_24222 ? T_47656_124 : GEN_2589;
  assign GEN_2591 = 9'h7d == T_24222 ? T_47656_125 : GEN_2590;
  assign GEN_2592 = 9'h7e == T_24222 ? T_47656_126 : GEN_2591;
  assign GEN_2593 = 9'h7f == T_24222 ? T_47656_127 : GEN_2592;
  assign GEN_2594 = 9'h80 == T_24222 ? T_47656_128 : GEN_2593;
  assign GEN_2595 = 9'h81 == T_24222 ? T_47656_129 : GEN_2594;
  assign GEN_2596 = 9'h82 == T_24222 ? T_47656_130 : GEN_2595;
  assign GEN_2597 = 9'h83 == T_24222 ? T_47656_131 : GEN_2596;
  assign GEN_2598 = 9'h84 == T_24222 ? T_47656_132 : GEN_2597;
  assign GEN_2599 = 9'h85 == T_24222 ? T_47656_133 : GEN_2598;
  assign GEN_2600 = 9'h86 == T_24222 ? T_47656_134 : GEN_2599;
  assign GEN_2601 = 9'h87 == T_24222 ? T_47656_135 : GEN_2600;
  assign GEN_2602 = 9'h88 == T_24222 ? T_47656_136 : GEN_2601;
  assign GEN_2603 = 9'h89 == T_24222 ? T_47656_137 : GEN_2602;
  assign GEN_2604 = 9'h8a == T_24222 ? T_47656_138 : GEN_2603;
  assign GEN_2605 = 9'h8b == T_24222 ? T_47656_139 : GEN_2604;
  assign GEN_2606 = 9'h8c == T_24222 ? T_47656_140 : GEN_2605;
  assign GEN_2607 = 9'h8d == T_24222 ? T_47656_141 : GEN_2606;
  assign GEN_2608 = 9'h8e == T_24222 ? T_47656_142 : GEN_2607;
  assign GEN_2609 = 9'h8f == T_24222 ? T_47656_143 : GEN_2608;
  assign GEN_2610 = 9'h90 == T_24222 ? T_47656_144 : GEN_2609;
  assign GEN_2611 = 9'h91 == T_24222 ? T_47656_145 : GEN_2610;
  assign GEN_2612 = 9'h92 == T_24222 ? T_47656_146 : GEN_2611;
  assign GEN_2613 = 9'h93 == T_24222 ? T_47656_147 : GEN_2612;
  assign GEN_2614 = 9'h94 == T_24222 ? T_47656_148 : GEN_2613;
  assign GEN_2615 = 9'h95 == T_24222 ? T_47656_149 : GEN_2614;
  assign GEN_2616 = 9'h96 == T_24222 ? T_47656_150 : GEN_2615;
  assign GEN_2617 = 9'h97 == T_24222 ? T_47656_151 : GEN_2616;
  assign GEN_2618 = 9'h98 == T_24222 ? T_47656_152 : GEN_2617;
  assign GEN_2619 = 9'h99 == T_24222 ? T_47656_153 : GEN_2618;
  assign GEN_2620 = 9'h9a == T_24222 ? T_47656_154 : GEN_2619;
  assign GEN_2621 = 9'h9b == T_24222 ? T_47656_155 : GEN_2620;
  assign GEN_2622 = 9'h9c == T_24222 ? T_47656_156 : GEN_2621;
  assign GEN_2623 = 9'h9d == T_24222 ? T_47656_157 : GEN_2622;
  assign GEN_2624 = 9'h9e == T_24222 ? T_47656_158 : GEN_2623;
  assign GEN_2625 = 9'h9f == T_24222 ? T_47656_159 : GEN_2624;
  assign GEN_2626 = 9'ha0 == T_24222 ? T_47656_160 : GEN_2625;
  assign GEN_2627 = 9'ha1 == T_24222 ? T_47656_161 : GEN_2626;
  assign GEN_2628 = 9'ha2 == T_24222 ? T_47656_162 : GEN_2627;
  assign GEN_2629 = 9'ha3 == T_24222 ? T_47656_163 : GEN_2628;
  assign GEN_2630 = 9'ha4 == T_24222 ? T_47656_164 : GEN_2629;
  assign GEN_2631 = 9'ha5 == T_24222 ? T_47656_165 : GEN_2630;
  assign GEN_2632 = 9'ha6 == T_24222 ? T_47656_166 : GEN_2631;
  assign GEN_2633 = 9'ha7 == T_24222 ? T_47656_167 : GEN_2632;
  assign GEN_2634 = 9'ha8 == T_24222 ? T_47656_168 : GEN_2633;
  assign GEN_2635 = 9'ha9 == T_24222 ? T_47656_169 : GEN_2634;
  assign GEN_2636 = 9'haa == T_24222 ? T_47656_170 : GEN_2635;
  assign GEN_2637 = 9'hab == T_24222 ? T_47656_171 : GEN_2636;
  assign GEN_2638 = 9'hac == T_24222 ? T_47656_172 : GEN_2637;
  assign GEN_2639 = 9'had == T_24222 ? T_47656_173 : GEN_2638;
  assign GEN_2640 = 9'hae == T_24222 ? T_47656_174 : GEN_2639;
  assign GEN_2641 = 9'haf == T_24222 ? T_47656_175 : GEN_2640;
  assign GEN_2642 = 9'hb0 == T_24222 ? T_47656_176 : GEN_2641;
  assign GEN_2643 = 9'hb1 == T_24222 ? T_47656_177 : GEN_2642;
  assign GEN_2644 = 9'hb2 == T_24222 ? T_47656_178 : GEN_2643;
  assign GEN_2645 = 9'hb3 == T_24222 ? T_47656_179 : GEN_2644;
  assign GEN_2646 = 9'hb4 == T_24222 ? T_47656_180 : GEN_2645;
  assign GEN_2647 = 9'hb5 == T_24222 ? T_47656_181 : GEN_2646;
  assign GEN_2648 = 9'hb6 == T_24222 ? T_47656_182 : GEN_2647;
  assign GEN_2649 = 9'hb7 == T_24222 ? T_47656_183 : GEN_2648;
  assign GEN_2650 = 9'hb8 == T_24222 ? T_47656_184 : GEN_2649;
  assign GEN_2651 = 9'hb9 == T_24222 ? T_47656_185 : GEN_2650;
  assign GEN_2652 = 9'hba == T_24222 ? T_47656_186 : GEN_2651;
  assign GEN_2653 = 9'hbb == T_24222 ? T_47656_187 : GEN_2652;
  assign GEN_2654 = 9'hbc == T_24222 ? T_47656_188 : GEN_2653;
  assign GEN_2655 = 9'hbd == T_24222 ? T_47656_189 : GEN_2654;
  assign GEN_2656 = 9'hbe == T_24222 ? T_47656_190 : GEN_2655;
  assign GEN_2657 = 9'hbf == T_24222 ? T_47656_191 : GEN_2656;
  assign GEN_2658 = 9'hc0 == T_24222 ? T_47656_192 : GEN_2657;
  assign GEN_2659 = 9'hc1 == T_24222 ? T_47656_193 : GEN_2658;
  assign GEN_2660 = 9'hc2 == T_24222 ? T_47656_194 : GEN_2659;
  assign GEN_2661 = 9'hc3 == T_24222 ? T_47656_195 : GEN_2660;
  assign GEN_2662 = 9'hc4 == T_24222 ? T_47656_196 : GEN_2661;
  assign GEN_2663 = 9'hc5 == T_24222 ? T_47656_197 : GEN_2662;
  assign GEN_2664 = 9'hc6 == T_24222 ? T_47656_198 : GEN_2663;
  assign GEN_2665 = 9'hc7 == T_24222 ? T_47656_199 : GEN_2664;
  assign GEN_2666 = 9'hc8 == T_24222 ? T_47656_200 : GEN_2665;
  assign GEN_2667 = 9'hc9 == T_24222 ? T_47656_201 : GEN_2666;
  assign GEN_2668 = 9'hca == T_24222 ? T_47656_202 : GEN_2667;
  assign GEN_2669 = 9'hcb == T_24222 ? T_47656_203 : GEN_2668;
  assign GEN_2670 = 9'hcc == T_24222 ? T_47656_204 : GEN_2669;
  assign GEN_2671 = 9'hcd == T_24222 ? T_47656_205 : GEN_2670;
  assign GEN_2672 = 9'hce == T_24222 ? T_47656_206 : GEN_2671;
  assign GEN_2673 = 9'hcf == T_24222 ? T_47656_207 : GEN_2672;
  assign GEN_2674 = 9'hd0 == T_24222 ? T_47656_208 : GEN_2673;
  assign GEN_2675 = 9'hd1 == T_24222 ? T_47656_209 : GEN_2674;
  assign GEN_2676 = 9'hd2 == T_24222 ? T_47656_210 : GEN_2675;
  assign GEN_2677 = 9'hd3 == T_24222 ? T_47656_211 : GEN_2676;
  assign GEN_2678 = 9'hd4 == T_24222 ? T_47656_212 : GEN_2677;
  assign GEN_2679 = 9'hd5 == T_24222 ? T_47656_213 : GEN_2678;
  assign GEN_2680 = 9'hd6 == T_24222 ? T_47656_214 : GEN_2679;
  assign GEN_2681 = 9'hd7 == T_24222 ? T_47656_215 : GEN_2680;
  assign GEN_2682 = 9'hd8 == T_24222 ? T_47656_216 : GEN_2681;
  assign GEN_2683 = 9'hd9 == T_24222 ? T_47656_217 : GEN_2682;
  assign GEN_2684 = 9'hda == T_24222 ? T_47656_218 : GEN_2683;
  assign GEN_2685 = 9'hdb == T_24222 ? T_47656_219 : GEN_2684;
  assign GEN_2686 = 9'hdc == T_24222 ? T_47656_220 : GEN_2685;
  assign GEN_2687 = 9'hdd == T_24222 ? T_47656_221 : GEN_2686;
  assign GEN_2688 = 9'hde == T_24222 ? T_47656_222 : GEN_2687;
  assign GEN_2689 = 9'hdf == T_24222 ? T_47656_223 : GEN_2688;
  assign GEN_2690 = 9'he0 == T_24222 ? T_47656_224 : GEN_2689;
  assign GEN_2691 = 9'he1 == T_24222 ? T_47656_225 : GEN_2690;
  assign GEN_2692 = 9'he2 == T_24222 ? T_47656_226 : GEN_2691;
  assign GEN_2693 = 9'he3 == T_24222 ? T_47656_227 : GEN_2692;
  assign GEN_2694 = 9'he4 == T_24222 ? T_47656_228 : GEN_2693;
  assign GEN_2695 = 9'he5 == T_24222 ? T_47656_229 : GEN_2694;
  assign GEN_2696 = 9'he6 == T_24222 ? T_47656_230 : GEN_2695;
  assign GEN_2697 = 9'he7 == T_24222 ? T_47656_231 : GEN_2696;
  assign GEN_2698 = 9'he8 == T_24222 ? T_47656_232 : GEN_2697;
  assign GEN_2699 = 9'he9 == T_24222 ? T_47656_233 : GEN_2698;
  assign GEN_2700 = 9'hea == T_24222 ? T_47656_234 : GEN_2699;
  assign GEN_2701 = 9'heb == T_24222 ? T_47656_235 : GEN_2700;
  assign GEN_2702 = 9'hec == T_24222 ? T_47656_236 : GEN_2701;
  assign GEN_2703 = 9'hed == T_24222 ? T_47656_237 : GEN_2702;
  assign GEN_2704 = 9'hee == T_24222 ? T_47656_238 : GEN_2703;
  assign GEN_2705 = 9'hef == T_24222 ? T_47656_239 : GEN_2704;
  assign GEN_2706 = 9'hf0 == T_24222 ? T_47656_240 : GEN_2705;
  assign GEN_2707 = 9'hf1 == T_24222 ? T_47656_241 : GEN_2706;
  assign GEN_2708 = 9'hf2 == T_24222 ? T_47656_242 : GEN_2707;
  assign GEN_2709 = 9'hf3 == T_24222 ? T_47656_243 : GEN_2708;
  assign GEN_2710 = 9'hf4 == T_24222 ? T_47656_244 : GEN_2709;
  assign GEN_2711 = 9'hf5 == T_24222 ? T_47656_245 : GEN_2710;
  assign GEN_2712 = 9'hf6 == T_24222 ? T_47656_246 : GEN_2711;
  assign GEN_2713 = 9'hf7 == T_24222 ? T_47656_247 : GEN_2712;
  assign GEN_2714 = 9'hf8 == T_24222 ? T_47656_248 : GEN_2713;
  assign GEN_2715 = 9'hf9 == T_24222 ? T_47656_249 : GEN_2714;
  assign GEN_2716 = 9'hfa == T_24222 ? T_47656_250 : GEN_2715;
  assign GEN_2717 = 9'hfb == T_24222 ? T_47656_251 : GEN_2716;
  assign GEN_2718 = 9'hfc == T_24222 ? T_47656_252 : GEN_2717;
  assign GEN_2719 = 9'hfd == T_24222 ? T_47656_253 : GEN_2718;
  assign GEN_2720 = 9'hfe == T_24222 ? T_47656_254 : GEN_2719;
  assign GEN_2721 = 9'hff == T_24222 ? T_47656_255 : GEN_2720;
  assign GEN_2722 = 9'h100 == T_24222 ? T_47656_256 : GEN_2721;
  assign GEN_2723 = 9'h101 == T_24222 ? T_47656_257 : GEN_2722;
  assign GEN_2724 = 9'h102 == T_24222 ? T_47656_258 : GEN_2723;
  assign GEN_2725 = 9'h103 == T_24222 ? T_47656_259 : GEN_2724;
  assign GEN_2726 = 9'h104 == T_24222 ? T_47656_260 : GEN_2725;
  assign GEN_2727 = 9'h105 == T_24222 ? T_47656_261 : GEN_2726;
  assign GEN_2728 = 9'h106 == T_24222 ? T_47656_262 : GEN_2727;
  assign GEN_2729 = 9'h107 == T_24222 ? T_47656_263 : GEN_2728;
  assign GEN_2730 = 9'h108 == T_24222 ? T_47656_264 : GEN_2729;
  assign GEN_2731 = 9'h109 == T_24222 ? T_47656_265 : GEN_2730;
  assign GEN_2732 = 9'h10a == T_24222 ? T_47656_266 : GEN_2731;
  assign GEN_2733 = 9'h10b == T_24222 ? T_47656_267 : GEN_2732;
  assign GEN_2734 = 9'h10c == T_24222 ? T_47656_268 : GEN_2733;
  assign GEN_2735 = 9'h10d == T_24222 ? T_47656_269 : GEN_2734;
  assign GEN_2736 = 9'h10e == T_24222 ? T_47656_270 : GEN_2735;
  assign GEN_2737 = 9'h10f == T_24222 ? T_47656_271 : GEN_2736;
  assign GEN_2738 = 9'h110 == T_24222 ? T_47656_272 : GEN_2737;
  assign GEN_2739 = 9'h111 == T_24222 ? T_47656_273 : GEN_2738;
  assign GEN_2740 = 9'h112 == T_24222 ? T_47656_274 : GEN_2739;
  assign GEN_2741 = 9'h113 == T_24222 ? T_47656_275 : GEN_2740;
  assign GEN_2742 = 9'h114 == T_24222 ? T_47656_276 : GEN_2741;
  assign GEN_2743 = 9'h115 == T_24222 ? T_47656_277 : GEN_2742;
  assign GEN_2744 = 9'h116 == T_24222 ? T_47656_278 : GEN_2743;
  assign GEN_2745 = 9'h117 == T_24222 ? T_47656_279 : GEN_2744;
  assign GEN_2746 = 9'h118 == T_24222 ? T_47656_280 : GEN_2745;
  assign GEN_2747 = 9'h119 == T_24222 ? T_47656_281 : GEN_2746;
  assign GEN_2748 = 9'h11a == T_24222 ? T_47656_282 : GEN_2747;
  assign GEN_2749 = 9'h11b == T_24222 ? T_47656_283 : GEN_2748;
  assign GEN_2750 = 9'h11c == T_24222 ? T_47656_284 : GEN_2749;
  assign GEN_2751 = 9'h11d == T_24222 ? T_47656_285 : GEN_2750;
  assign GEN_2752 = 9'h11e == T_24222 ? T_47656_286 : GEN_2751;
  assign GEN_2753 = 9'h11f == T_24222 ? T_47656_287 : GEN_2752;
  assign GEN_2754 = 9'h120 == T_24222 ? T_47656_288 : GEN_2753;
  assign GEN_2755 = 9'h121 == T_24222 ? T_47656_289 : GEN_2754;
  assign GEN_2756 = 9'h122 == T_24222 ? T_47656_290 : GEN_2755;
  assign GEN_2757 = 9'h123 == T_24222 ? T_47656_291 : GEN_2756;
  assign GEN_2758 = 9'h124 == T_24222 ? T_47656_292 : GEN_2757;
  assign GEN_2759 = 9'h125 == T_24222 ? T_47656_293 : GEN_2758;
  assign GEN_2760 = 9'h126 == T_24222 ? T_47656_294 : GEN_2759;
  assign GEN_2761 = 9'h127 == T_24222 ? T_47656_295 : GEN_2760;
  assign GEN_2762 = 9'h128 == T_24222 ? T_47656_296 : GEN_2761;
  assign GEN_2763 = 9'h129 == T_24222 ? T_47656_297 : GEN_2762;
  assign GEN_2764 = 9'h12a == T_24222 ? T_47656_298 : GEN_2763;
  assign GEN_2765 = 9'h12b == T_24222 ? T_47656_299 : GEN_2764;
  assign GEN_2766 = 9'h12c == T_24222 ? T_47656_300 : GEN_2765;
  assign GEN_2767 = 9'h12d == T_24222 ? T_47656_301 : GEN_2766;
  assign GEN_2768 = 9'h12e == T_24222 ? T_47656_302 : GEN_2767;
  assign GEN_2769 = 9'h12f == T_24222 ? T_47656_303 : GEN_2768;
  assign GEN_2770 = 9'h130 == T_24222 ? T_47656_304 : GEN_2769;
  assign GEN_2771 = 9'h131 == T_24222 ? T_47656_305 : GEN_2770;
  assign GEN_2772 = 9'h132 == T_24222 ? T_47656_306 : GEN_2771;
  assign GEN_2773 = 9'h133 == T_24222 ? T_47656_307 : GEN_2772;
  assign GEN_2774 = 9'h134 == T_24222 ? T_47656_308 : GEN_2773;
  assign GEN_2775 = 9'h135 == T_24222 ? T_47656_309 : GEN_2774;
  assign GEN_2776 = 9'h136 == T_24222 ? T_47656_310 : GEN_2775;
  assign GEN_2777 = 9'h137 == T_24222 ? T_47656_311 : GEN_2776;
  assign GEN_2778 = 9'h138 == T_24222 ? T_47656_312 : GEN_2777;
  assign GEN_2779 = 9'h139 == T_24222 ? T_47656_313 : GEN_2778;
  assign GEN_2780 = 9'h13a == T_24222 ? T_47656_314 : GEN_2779;
  assign GEN_2781 = 9'h13b == T_24222 ? T_47656_315 : GEN_2780;
  assign GEN_2782 = 9'h13c == T_24222 ? T_47656_316 : GEN_2781;
  assign GEN_2783 = 9'h13d == T_24222 ? T_47656_317 : GEN_2782;
  assign GEN_2784 = 9'h13e == T_24222 ? T_47656_318 : GEN_2783;
  assign GEN_2785 = 9'h13f == T_24222 ? T_47656_319 : GEN_2784;
  assign GEN_2786 = 9'h140 == T_24222 ? T_47656_320 : GEN_2785;
  assign GEN_2787 = 9'h141 == T_24222 ? T_47656_321 : GEN_2786;
  assign GEN_2788 = 9'h142 == T_24222 ? T_47656_322 : GEN_2787;
  assign GEN_2789 = 9'h143 == T_24222 ? T_47656_323 : GEN_2788;
  assign GEN_2790 = 9'h144 == T_24222 ? T_47656_324 : GEN_2789;
  assign GEN_2791 = 9'h145 == T_24222 ? T_47656_325 : GEN_2790;
  assign GEN_2792 = 9'h146 == T_24222 ? T_47656_326 : GEN_2791;
  assign GEN_2793 = 9'h147 == T_24222 ? T_47656_327 : GEN_2792;
  assign GEN_2794 = 9'h148 == T_24222 ? T_47656_328 : GEN_2793;
  assign GEN_2795 = 9'h149 == T_24222 ? T_47656_329 : GEN_2794;
  assign GEN_2796 = 9'h14a == T_24222 ? T_47656_330 : GEN_2795;
  assign GEN_2797 = 9'h14b == T_24222 ? T_47656_331 : GEN_2796;
  assign GEN_2798 = 9'h14c == T_24222 ? T_47656_332 : GEN_2797;
  assign GEN_2799 = 9'h14d == T_24222 ? T_47656_333 : GEN_2798;
  assign GEN_2800 = 9'h14e == T_24222 ? T_47656_334 : GEN_2799;
  assign GEN_2801 = 9'h14f == T_24222 ? T_47656_335 : GEN_2800;
  assign GEN_2802 = 9'h150 == T_24222 ? T_47656_336 : GEN_2801;
  assign GEN_2803 = 9'h151 == T_24222 ? T_47656_337 : GEN_2802;
  assign GEN_2804 = 9'h152 == T_24222 ? T_47656_338 : GEN_2803;
  assign GEN_2805 = 9'h153 == T_24222 ? T_47656_339 : GEN_2804;
  assign GEN_2806 = 9'h154 == T_24222 ? T_47656_340 : GEN_2805;
  assign GEN_2807 = 9'h155 == T_24222 ? T_47656_341 : GEN_2806;
  assign GEN_2808 = 9'h156 == T_24222 ? T_47656_342 : GEN_2807;
  assign GEN_2809 = 9'h157 == T_24222 ? T_47656_343 : GEN_2808;
  assign GEN_2810 = 9'h158 == T_24222 ? T_47656_344 : GEN_2809;
  assign GEN_2811 = 9'h159 == T_24222 ? T_47656_345 : GEN_2810;
  assign GEN_2812 = 9'h15a == T_24222 ? T_47656_346 : GEN_2811;
  assign GEN_2813 = 9'h15b == T_24222 ? T_47656_347 : GEN_2812;
  assign GEN_2814 = 9'h15c == T_24222 ? T_47656_348 : GEN_2813;
  assign GEN_2815 = 9'h15d == T_24222 ? T_47656_349 : GEN_2814;
  assign GEN_2816 = 9'h15e == T_24222 ? T_47656_350 : GEN_2815;
  assign GEN_2817 = 9'h15f == T_24222 ? T_47656_351 : GEN_2816;
  assign GEN_2818 = 9'h160 == T_24222 ? T_47656_352 : GEN_2817;
  assign GEN_2819 = 9'h161 == T_24222 ? T_47656_353 : GEN_2818;
  assign GEN_2820 = 9'h162 == T_24222 ? T_47656_354 : GEN_2819;
  assign GEN_2821 = 9'h163 == T_24222 ? T_47656_355 : GEN_2820;
  assign GEN_2822 = 9'h164 == T_24222 ? T_47656_356 : GEN_2821;
  assign GEN_2823 = 9'h165 == T_24222 ? T_47656_357 : GEN_2822;
  assign GEN_2824 = 9'h166 == T_24222 ? T_47656_358 : GEN_2823;
  assign GEN_2825 = 9'h167 == T_24222 ? T_47656_359 : GEN_2824;
  assign GEN_2826 = 9'h168 == T_24222 ? T_47656_360 : GEN_2825;
  assign GEN_2827 = 9'h169 == T_24222 ? T_47656_361 : GEN_2826;
  assign GEN_2828 = 9'h16a == T_24222 ? T_47656_362 : GEN_2827;
  assign GEN_2829 = 9'h16b == T_24222 ? T_47656_363 : GEN_2828;
  assign GEN_2830 = 9'h16c == T_24222 ? T_47656_364 : GEN_2829;
  assign GEN_2831 = 9'h16d == T_24222 ? T_47656_365 : GEN_2830;
  assign GEN_2832 = 9'h16e == T_24222 ? T_47656_366 : GEN_2831;
  assign GEN_2833 = 9'h16f == T_24222 ? T_47656_367 : GEN_2832;
  assign GEN_2834 = 9'h170 == T_24222 ? T_47656_368 : GEN_2833;
  assign GEN_2835 = 9'h171 == T_24222 ? T_47656_369 : GEN_2834;
  assign GEN_2836 = 9'h172 == T_24222 ? T_47656_370 : GEN_2835;
  assign GEN_2837 = 9'h173 == T_24222 ? T_47656_371 : GEN_2836;
  assign GEN_2838 = 9'h174 == T_24222 ? T_47656_372 : GEN_2837;
  assign GEN_2839 = 9'h175 == T_24222 ? T_47656_373 : GEN_2838;
  assign GEN_2840 = 9'h176 == T_24222 ? T_47656_374 : GEN_2839;
  assign GEN_2841 = 9'h177 == T_24222 ? T_47656_375 : GEN_2840;
  assign GEN_2842 = 9'h178 == T_24222 ? T_47656_376 : GEN_2841;
  assign GEN_2843 = 9'h179 == T_24222 ? T_47656_377 : GEN_2842;
  assign GEN_2844 = 9'h17a == T_24222 ? T_47656_378 : GEN_2843;
  assign GEN_2845 = 9'h17b == T_24222 ? T_47656_379 : GEN_2844;
  assign GEN_2846 = 9'h17c == T_24222 ? T_47656_380 : GEN_2845;
  assign GEN_2847 = 9'h17d == T_24222 ? T_47656_381 : GEN_2846;
  assign GEN_2848 = 9'h17e == T_24222 ? T_47656_382 : GEN_2847;
  assign GEN_2849 = 9'h17f == T_24222 ? T_47656_383 : GEN_2848;
  assign GEN_2850 = 9'h180 == T_24222 ? T_47656_384 : GEN_2849;
  assign GEN_2851 = 9'h181 == T_24222 ? T_47656_385 : GEN_2850;
  assign GEN_2852 = 9'h182 == T_24222 ? T_47656_386 : GEN_2851;
  assign GEN_2853 = 9'h183 == T_24222 ? T_47656_387 : GEN_2852;
  assign GEN_2854 = 9'h184 == T_24222 ? T_47656_388 : GEN_2853;
  assign GEN_2855 = 9'h185 == T_24222 ? T_47656_389 : GEN_2854;
  assign GEN_2856 = 9'h186 == T_24222 ? T_47656_390 : GEN_2855;
  assign GEN_2857 = 9'h187 == T_24222 ? T_47656_391 : GEN_2856;
  assign GEN_2858 = 9'h188 == T_24222 ? T_47656_392 : GEN_2857;
  assign GEN_2859 = 9'h189 == T_24222 ? T_47656_393 : GEN_2858;
  assign GEN_2860 = 9'h18a == T_24222 ? T_47656_394 : GEN_2859;
  assign GEN_2861 = 9'h18b == T_24222 ? T_47656_395 : GEN_2860;
  assign GEN_2862 = 9'h18c == T_24222 ? T_47656_396 : GEN_2861;
  assign GEN_2863 = 9'h18d == T_24222 ? T_47656_397 : GEN_2862;
  assign GEN_2864 = 9'h18e == T_24222 ? T_47656_398 : GEN_2863;
  assign GEN_2865 = 9'h18f == T_24222 ? T_47656_399 : GEN_2864;
  assign GEN_2866 = 9'h190 == T_24222 ? T_47656_400 : GEN_2865;
  assign GEN_2867 = 9'h191 == T_24222 ? T_47656_401 : GEN_2866;
  assign GEN_2868 = 9'h192 == T_24222 ? T_47656_402 : GEN_2867;
  assign GEN_2869 = 9'h193 == T_24222 ? T_47656_403 : GEN_2868;
  assign GEN_2870 = 9'h194 == T_24222 ? T_47656_404 : GEN_2869;
  assign GEN_2871 = 9'h195 == T_24222 ? T_47656_405 : GEN_2870;
  assign GEN_2872 = 9'h196 == T_24222 ? T_47656_406 : GEN_2871;
  assign GEN_2873 = 9'h197 == T_24222 ? T_47656_407 : GEN_2872;
  assign GEN_2874 = 9'h198 == T_24222 ? T_47656_408 : GEN_2873;
  assign GEN_2875 = 9'h199 == T_24222 ? T_47656_409 : GEN_2874;
  assign GEN_2876 = 9'h19a == T_24222 ? T_47656_410 : GEN_2875;
  assign GEN_2877 = 9'h19b == T_24222 ? T_47656_411 : GEN_2876;
  assign GEN_2878 = 9'h19c == T_24222 ? T_47656_412 : GEN_2877;
  assign GEN_2879 = 9'h19d == T_24222 ? T_47656_413 : GEN_2878;
  assign GEN_2880 = 9'h19e == T_24222 ? T_47656_414 : GEN_2879;
  assign GEN_2881 = 9'h19f == T_24222 ? T_47656_415 : GEN_2880;
  assign GEN_2882 = 9'h1a0 == T_24222 ? T_47656_416 : GEN_2881;
  assign GEN_2883 = 9'h1a1 == T_24222 ? T_47656_417 : GEN_2882;
  assign GEN_2884 = 9'h1a2 == T_24222 ? T_47656_418 : GEN_2883;
  assign GEN_2885 = 9'h1a3 == T_24222 ? T_47656_419 : GEN_2884;
  assign GEN_2886 = 9'h1a4 == T_24222 ? T_47656_420 : GEN_2885;
  assign GEN_2887 = 9'h1a5 == T_24222 ? T_47656_421 : GEN_2886;
  assign GEN_2888 = 9'h1a6 == T_24222 ? T_47656_422 : GEN_2887;
  assign GEN_2889 = 9'h1a7 == T_24222 ? T_47656_423 : GEN_2888;
  assign GEN_2890 = 9'h1a8 == T_24222 ? T_47656_424 : GEN_2889;
  assign GEN_2891 = 9'h1a9 == T_24222 ? T_47656_425 : GEN_2890;
  assign GEN_2892 = 9'h1aa == T_24222 ? T_47656_426 : GEN_2891;
  assign GEN_2893 = 9'h1ab == T_24222 ? T_47656_427 : GEN_2892;
  assign GEN_2894 = 9'h1ac == T_24222 ? T_47656_428 : GEN_2893;
  assign GEN_2895 = 9'h1ad == T_24222 ? T_47656_429 : GEN_2894;
  assign GEN_2896 = 9'h1ae == T_24222 ? T_47656_430 : GEN_2895;
  assign GEN_2897 = 9'h1af == T_24222 ? T_47656_431 : GEN_2896;
  assign GEN_2898 = 9'h1b0 == T_24222 ? T_47656_432 : GEN_2897;
  assign GEN_2899 = 9'h1b1 == T_24222 ? T_47656_433 : GEN_2898;
  assign GEN_2900 = 9'h1b2 == T_24222 ? T_47656_434 : GEN_2899;
  assign GEN_2901 = 9'h1b3 == T_24222 ? T_47656_435 : GEN_2900;
  assign GEN_2902 = 9'h1b4 == T_24222 ? T_47656_436 : GEN_2901;
  assign GEN_2903 = 9'h1b5 == T_24222 ? T_47656_437 : GEN_2902;
  assign GEN_2904 = 9'h1b6 == T_24222 ? T_47656_438 : GEN_2903;
  assign GEN_2905 = 9'h1b7 == T_24222 ? T_47656_439 : GEN_2904;
  assign GEN_2906 = 9'h1b8 == T_24222 ? T_47656_440 : GEN_2905;
  assign GEN_2907 = 9'h1b9 == T_24222 ? T_47656_441 : GEN_2906;
  assign GEN_2908 = 9'h1ba == T_24222 ? T_47656_442 : GEN_2907;
  assign GEN_2909 = 9'h1bb == T_24222 ? T_47656_443 : GEN_2908;
  assign GEN_2910 = 9'h1bc == T_24222 ? T_47656_444 : GEN_2909;
  assign GEN_2911 = 9'h1bd == T_24222 ? T_47656_445 : GEN_2910;
  assign GEN_2912 = 9'h1be == T_24222 ? T_47656_446 : GEN_2911;
  assign GEN_2913 = 9'h1bf == T_24222 ? T_47656_447 : GEN_2912;
  assign GEN_2914 = 9'h1c0 == T_24222 ? T_47656_448 : GEN_2913;
  assign GEN_2915 = 9'h1c1 == T_24222 ? T_47656_449 : GEN_2914;
  assign GEN_2916 = 9'h1c2 == T_24222 ? T_47656_450 : GEN_2915;
  assign GEN_2917 = 9'h1c3 == T_24222 ? T_47656_451 : GEN_2916;
  assign GEN_2918 = 9'h1c4 == T_24222 ? T_47656_452 : GEN_2917;
  assign GEN_2919 = 9'h1c5 == T_24222 ? T_47656_453 : GEN_2918;
  assign GEN_2920 = 9'h1c6 == T_24222 ? T_47656_454 : GEN_2919;
  assign GEN_2921 = 9'h1c7 == T_24222 ? T_47656_455 : GEN_2920;
  assign GEN_2922 = 9'h1c8 == T_24222 ? T_47656_456 : GEN_2921;
  assign GEN_2923 = 9'h1c9 == T_24222 ? T_47656_457 : GEN_2922;
  assign GEN_2924 = 9'h1ca == T_24222 ? T_47656_458 : GEN_2923;
  assign GEN_2925 = 9'h1cb == T_24222 ? T_47656_459 : GEN_2924;
  assign GEN_2926 = 9'h1cc == T_24222 ? T_47656_460 : GEN_2925;
  assign GEN_2927 = 9'h1cd == T_24222 ? T_47656_461 : GEN_2926;
  assign GEN_2928 = 9'h1ce == T_24222 ? T_47656_462 : GEN_2927;
  assign GEN_2929 = 9'h1cf == T_24222 ? T_47656_463 : GEN_2928;
  assign GEN_2930 = 9'h1d0 == T_24222 ? T_47656_464 : GEN_2929;
  assign GEN_2931 = 9'h1d1 == T_24222 ? T_47656_465 : GEN_2930;
  assign GEN_2932 = 9'h1d2 == T_24222 ? T_47656_466 : GEN_2931;
  assign GEN_2933 = 9'h1d3 == T_24222 ? T_47656_467 : GEN_2932;
  assign GEN_2934 = 9'h1d4 == T_24222 ? T_47656_468 : GEN_2933;
  assign GEN_2935 = 9'h1d5 == T_24222 ? T_47656_469 : GEN_2934;
  assign GEN_2936 = 9'h1d6 == T_24222 ? T_47656_470 : GEN_2935;
  assign GEN_2937 = 9'h1d7 == T_24222 ? T_47656_471 : GEN_2936;
  assign GEN_2938 = 9'h1d8 == T_24222 ? T_47656_472 : GEN_2937;
  assign GEN_2939 = 9'h1d9 == T_24222 ? T_47656_473 : GEN_2938;
  assign GEN_2940 = 9'h1da == T_24222 ? T_47656_474 : GEN_2939;
  assign GEN_2941 = 9'h1db == T_24222 ? T_47656_475 : GEN_2940;
  assign GEN_2942 = 9'h1dc == T_24222 ? T_47656_476 : GEN_2941;
  assign GEN_2943 = 9'h1dd == T_24222 ? T_47656_477 : GEN_2942;
  assign GEN_2944 = 9'h1de == T_24222 ? T_47656_478 : GEN_2943;
  assign GEN_2945 = 9'h1df == T_24222 ? T_47656_479 : GEN_2944;
  assign GEN_2946 = 9'h1e0 == T_24222 ? T_47656_480 : GEN_2945;
  assign GEN_2947 = 9'h1e1 == T_24222 ? T_47656_481 : GEN_2946;
  assign GEN_2948 = 9'h1e2 == T_24222 ? T_47656_482 : GEN_2947;
  assign GEN_2949 = 9'h1e3 == T_24222 ? T_47656_483 : GEN_2948;
  assign GEN_2950 = 9'h1e4 == T_24222 ? T_47656_484 : GEN_2949;
  assign GEN_2951 = 9'h1e5 == T_24222 ? T_47656_485 : GEN_2950;
  assign GEN_2952 = 9'h1e6 == T_24222 ? T_47656_486 : GEN_2951;
  assign GEN_2953 = 9'h1e7 == T_24222 ? T_47656_487 : GEN_2952;
  assign GEN_2954 = 9'h1e8 == T_24222 ? T_47656_488 : GEN_2953;
  assign GEN_2955 = 9'h1e9 == T_24222 ? T_47656_489 : GEN_2954;
  assign GEN_2956 = 9'h1ea == T_24222 ? T_47656_490 : GEN_2955;
  assign GEN_2957 = 9'h1eb == T_24222 ? T_47656_491 : GEN_2956;
  assign GEN_2958 = 9'h1ec == T_24222 ? T_47656_492 : GEN_2957;
  assign GEN_2959 = 9'h1ed == T_24222 ? T_47656_493 : GEN_2958;
  assign GEN_2960 = 9'h1ee == T_24222 ? T_47656_494 : GEN_2959;
  assign GEN_2961 = 9'h1ef == T_24222 ? T_47656_495 : GEN_2960;
  assign GEN_2962 = 9'h1f0 == T_24222 ? T_47656_496 : GEN_2961;
  assign GEN_2963 = 9'h1f1 == T_24222 ? T_47656_497 : GEN_2962;
  assign GEN_2964 = 9'h1f2 == T_24222 ? T_47656_498 : GEN_2963;
  assign GEN_2965 = 9'h1f3 == T_24222 ? T_47656_499 : GEN_2964;
  assign GEN_2966 = 9'h1f4 == T_24222 ? T_47656_500 : GEN_2965;
  assign GEN_2967 = 9'h1f5 == T_24222 ? T_47656_501 : GEN_2966;
  assign GEN_2968 = 9'h1f6 == T_24222 ? T_47656_502 : GEN_2967;
  assign GEN_2969 = 9'h1f7 == T_24222 ? T_47656_503 : GEN_2968;
  assign GEN_2970 = 9'h1f8 == T_24222 ? T_47656_504 : GEN_2969;
  assign GEN_2971 = 9'h1f9 == T_24222 ? T_47656_505 : GEN_2970;
  assign GEN_2972 = 9'h1fa == T_24222 ? T_47656_506 : GEN_2971;
  assign GEN_2973 = 9'h1fb == T_24222 ? T_47656_507 : GEN_2972;
  assign GEN_2974 = 9'h1fc == T_24222 ? T_47656_508 : GEN_2973;
  assign GEN_2975 = 9'h1fd == T_24222 ? T_47656_509 : GEN_2974;
  assign GEN_2976 = 9'h1fe == T_24222 ? T_47656_510 : GEN_2975;
  assign GEN_2977 = 9'h1ff == T_24222 ? T_47656_511 : GEN_2976;
  assign GEN_8 = GEN_3488;
  assign GEN_2978 = 9'h1 == T_24222 ? T_48687_1 : T_48687_0;
  assign GEN_2979 = 9'h2 == T_24222 ? T_48687_2 : GEN_2978;
  assign GEN_2980 = 9'h3 == T_24222 ? T_48687_3 : GEN_2979;
  assign GEN_2981 = 9'h4 == T_24222 ? T_48687_4 : GEN_2980;
  assign GEN_2982 = 9'h5 == T_24222 ? T_48687_5 : GEN_2981;
  assign GEN_2983 = 9'h6 == T_24222 ? T_48687_6 : GEN_2982;
  assign GEN_2984 = 9'h7 == T_24222 ? T_48687_7 : GEN_2983;
  assign GEN_2985 = 9'h8 == T_24222 ? T_48687_8 : GEN_2984;
  assign GEN_2986 = 9'h9 == T_24222 ? T_48687_9 : GEN_2985;
  assign GEN_2987 = 9'ha == T_24222 ? T_48687_10 : GEN_2986;
  assign GEN_2988 = 9'hb == T_24222 ? T_48687_11 : GEN_2987;
  assign GEN_2989 = 9'hc == T_24222 ? T_48687_12 : GEN_2988;
  assign GEN_2990 = 9'hd == T_24222 ? T_48687_13 : GEN_2989;
  assign GEN_2991 = 9'he == T_24222 ? T_48687_14 : GEN_2990;
  assign GEN_2992 = 9'hf == T_24222 ? T_48687_15 : GEN_2991;
  assign GEN_2993 = 9'h10 == T_24222 ? T_48687_16 : GEN_2992;
  assign GEN_2994 = 9'h11 == T_24222 ? T_48687_17 : GEN_2993;
  assign GEN_2995 = 9'h12 == T_24222 ? T_48687_18 : GEN_2994;
  assign GEN_2996 = 9'h13 == T_24222 ? T_48687_19 : GEN_2995;
  assign GEN_2997 = 9'h14 == T_24222 ? T_48687_20 : GEN_2996;
  assign GEN_2998 = 9'h15 == T_24222 ? T_48687_21 : GEN_2997;
  assign GEN_2999 = 9'h16 == T_24222 ? T_48687_22 : GEN_2998;
  assign GEN_3000 = 9'h17 == T_24222 ? T_48687_23 : GEN_2999;
  assign GEN_3001 = 9'h18 == T_24222 ? T_48687_24 : GEN_3000;
  assign GEN_3002 = 9'h19 == T_24222 ? T_48687_25 : GEN_3001;
  assign GEN_3003 = 9'h1a == T_24222 ? T_48687_26 : GEN_3002;
  assign GEN_3004 = 9'h1b == T_24222 ? T_48687_27 : GEN_3003;
  assign GEN_3005 = 9'h1c == T_24222 ? T_48687_28 : GEN_3004;
  assign GEN_3006 = 9'h1d == T_24222 ? T_48687_29 : GEN_3005;
  assign GEN_3007 = 9'h1e == T_24222 ? T_48687_30 : GEN_3006;
  assign GEN_3008 = 9'h1f == T_24222 ? T_48687_31 : GEN_3007;
  assign GEN_3009 = 9'h20 == T_24222 ? T_48687_32 : GEN_3008;
  assign GEN_3010 = 9'h21 == T_24222 ? T_48687_33 : GEN_3009;
  assign GEN_3011 = 9'h22 == T_24222 ? T_48687_34 : GEN_3010;
  assign GEN_3012 = 9'h23 == T_24222 ? T_48687_35 : GEN_3011;
  assign GEN_3013 = 9'h24 == T_24222 ? T_48687_36 : GEN_3012;
  assign GEN_3014 = 9'h25 == T_24222 ? T_48687_37 : GEN_3013;
  assign GEN_3015 = 9'h26 == T_24222 ? T_48687_38 : GEN_3014;
  assign GEN_3016 = 9'h27 == T_24222 ? T_48687_39 : GEN_3015;
  assign GEN_3017 = 9'h28 == T_24222 ? T_48687_40 : GEN_3016;
  assign GEN_3018 = 9'h29 == T_24222 ? T_48687_41 : GEN_3017;
  assign GEN_3019 = 9'h2a == T_24222 ? T_48687_42 : GEN_3018;
  assign GEN_3020 = 9'h2b == T_24222 ? T_48687_43 : GEN_3019;
  assign GEN_3021 = 9'h2c == T_24222 ? T_48687_44 : GEN_3020;
  assign GEN_3022 = 9'h2d == T_24222 ? T_48687_45 : GEN_3021;
  assign GEN_3023 = 9'h2e == T_24222 ? T_48687_46 : GEN_3022;
  assign GEN_3024 = 9'h2f == T_24222 ? T_48687_47 : GEN_3023;
  assign GEN_3025 = 9'h30 == T_24222 ? T_48687_48 : GEN_3024;
  assign GEN_3026 = 9'h31 == T_24222 ? T_48687_49 : GEN_3025;
  assign GEN_3027 = 9'h32 == T_24222 ? T_48687_50 : GEN_3026;
  assign GEN_3028 = 9'h33 == T_24222 ? T_48687_51 : GEN_3027;
  assign GEN_3029 = 9'h34 == T_24222 ? T_48687_52 : GEN_3028;
  assign GEN_3030 = 9'h35 == T_24222 ? T_48687_53 : GEN_3029;
  assign GEN_3031 = 9'h36 == T_24222 ? T_48687_54 : GEN_3030;
  assign GEN_3032 = 9'h37 == T_24222 ? T_48687_55 : GEN_3031;
  assign GEN_3033 = 9'h38 == T_24222 ? T_48687_56 : GEN_3032;
  assign GEN_3034 = 9'h39 == T_24222 ? T_48687_57 : GEN_3033;
  assign GEN_3035 = 9'h3a == T_24222 ? T_48687_58 : GEN_3034;
  assign GEN_3036 = 9'h3b == T_24222 ? T_48687_59 : GEN_3035;
  assign GEN_3037 = 9'h3c == T_24222 ? T_48687_60 : GEN_3036;
  assign GEN_3038 = 9'h3d == T_24222 ? T_48687_61 : GEN_3037;
  assign GEN_3039 = 9'h3e == T_24222 ? T_48687_62 : GEN_3038;
  assign GEN_3040 = 9'h3f == T_24222 ? T_48687_63 : GEN_3039;
  assign GEN_3041 = 9'h40 == T_24222 ? T_48687_64 : GEN_3040;
  assign GEN_3042 = 9'h41 == T_24222 ? T_48687_65 : GEN_3041;
  assign GEN_3043 = 9'h42 == T_24222 ? T_48687_66 : GEN_3042;
  assign GEN_3044 = 9'h43 == T_24222 ? T_48687_67 : GEN_3043;
  assign GEN_3045 = 9'h44 == T_24222 ? T_48687_68 : GEN_3044;
  assign GEN_3046 = 9'h45 == T_24222 ? T_48687_69 : GEN_3045;
  assign GEN_3047 = 9'h46 == T_24222 ? T_48687_70 : GEN_3046;
  assign GEN_3048 = 9'h47 == T_24222 ? T_48687_71 : GEN_3047;
  assign GEN_3049 = 9'h48 == T_24222 ? T_48687_72 : GEN_3048;
  assign GEN_3050 = 9'h49 == T_24222 ? T_48687_73 : GEN_3049;
  assign GEN_3051 = 9'h4a == T_24222 ? T_48687_74 : GEN_3050;
  assign GEN_3052 = 9'h4b == T_24222 ? T_48687_75 : GEN_3051;
  assign GEN_3053 = 9'h4c == T_24222 ? T_48687_76 : GEN_3052;
  assign GEN_3054 = 9'h4d == T_24222 ? T_48687_77 : GEN_3053;
  assign GEN_3055 = 9'h4e == T_24222 ? T_48687_78 : GEN_3054;
  assign GEN_3056 = 9'h4f == T_24222 ? T_48687_79 : GEN_3055;
  assign GEN_3057 = 9'h50 == T_24222 ? T_48687_80 : GEN_3056;
  assign GEN_3058 = 9'h51 == T_24222 ? T_48687_81 : GEN_3057;
  assign GEN_3059 = 9'h52 == T_24222 ? T_48687_82 : GEN_3058;
  assign GEN_3060 = 9'h53 == T_24222 ? T_48687_83 : GEN_3059;
  assign GEN_3061 = 9'h54 == T_24222 ? T_48687_84 : GEN_3060;
  assign GEN_3062 = 9'h55 == T_24222 ? T_48687_85 : GEN_3061;
  assign GEN_3063 = 9'h56 == T_24222 ? T_48687_86 : GEN_3062;
  assign GEN_3064 = 9'h57 == T_24222 ? T_48687_87 : GEN_3063;
  assign GEN_3065 = 9'h58 == T_24222 ? T_48687_88 : GEN_3064;
  assign GEN_3066 = 9'h59 == T_24222 ? T_48687_89 : GEN_3065;
  assign GEN_3067 = 9'h5a == T_24222 ? T_48687_90 : GEN_3066;
  assign GEN_3068 = 9'h5b == T_24222 ? T_48687_91 : GEN_3067;
  assign GEN_3069 = 9'h5c == T_24222 ? T_48687_92 : GEN_3068;
  assign GEN_3070 = 9'h5d == T_24222 ? T_48687_93 : GEN_3069;
  assign GEN_3071 = 9'h5e == T_24222 ? T_48687_94 : GEN_3070;
  assign GEN_3072 = 9'h5f == T_24222 ? T_48687_95 : GEN_3071;
  assign GEN_3073 = 9'h60 == T_24222 ? T_48687_96 : GEN_3072;
  assign GEN_3074 = 9'h61 == T_24222 ? T_48687_97 : GEN_3073;
  assign GEN_3075 = 9'h62 == T_24222 ? T_48687_98 : GEN_3074;
  assign GEN_3076 = 9'h63 == T_24222 ? T_48687_99 : GEN_3075;
  assign GEN_3077 = 9'h64 == T_24222 ? T_48687_100 : GEN_3076;
  assign GEN_3078 = 9'h65 == T_24222 ? T_48687_101 : GEN_3077;
  assign GEN_3079 = 9'h66 == T_24222 ? T_48687_102 : GEN_3078;
  assign GEN_3080 = 9'h67 == T_24222 ? T_48687_103 : GEN_3079;
  assign GEN_3081 = 9'h68 == T_24222 ? T_48687_104 : GEN_3080;
  assign GEN_3082 = 9'h69 == T_24222 ? T_48687_105 : GEN_3081;
  assign GEN_3083 = 9'h6a == T_24222 ? T_48687_106 : GEN_3082;
  assign GEN_3084 = 9'h6b == T_24222 ? T_48687_107 : GEN_3083;
  assign GEN_3085 = 9'h6c == T_24222 ? T_48687_108 : GEN_3084;
  assign GEN_3086 = 9'h6d == T_24222 ? T_48687_109 : GEN_3085;
  assign GEN_3087 = 9'h6e == T_24222 ? T_48687_110 : GEN_3086;
  assign GEN_3088 = 9'h6f == T_24222 ? T_48687_111 : GEN_3087;
  assign GEN_3089 = 9'h70 == T_24222 ? T_48687_112 : GEN_3088;
  assign GEN_3090 = 9'h71 == T_24222 ? T_48687_113 : GEN_3089;
  assign GEN_3091 = 9'h72 == T_24222 ? T_48687_114 : GEN_3090;
  assign GEN_3092 = 9'h73 == T_24222 ? T_48687_115 : GEN_3091;
  assign GEN_3093 = 9'h74 == T_24222 ? T_48687_116 : GEN_3092;
  assign GEN_3094 = 9'h75 == T_24222 ? T_48687_117 : GEN_3093;
  assign GEN_3095 = 9'h76 == T_24222 ? T_48687_118 : GEN_3094;
  assign GEN_3096 = 9'h77 == T_24222 ? T_48687_119 : GEN_3095;
  assign GEN_3097 = 9'h78 == T_24222 ? T_48687_120 : GEN_3096;
  assign GEN_3098 = 9'h79 == T_24222 ? T_48687_121 : GEN_3097;
  assign GEN_3099 = 9'h7a == T_24222 ? T_48687_122 : GEN_3098;
  assign GEN_3100 = 9'h7b == T_24222 ? T_48687_123 : GEN_3099;
  assign GEN_3101 = 9'h7c == T_24222 ? T_48687_124 : GEN_3100;
  assign GEN_3102 = 9'h7d == T_24222 ? T_48687_125 : GEN_3101;
  assign GEN_3103 = 9'h7e == T_24222 ? T_48687_126 : GEN_3102;
  assign GEN_3104 = 9'h7f == T_24222 ? T_48687_127 : GEN_3103;
  assign GEN_3105 = 9'h80 == T_24222 ? T_48687_128 : GEN_3104;
  assign GEN_3106 = 9'h81 == T_24222 ? T_48687_129 : GEN_3105;
  assign GEN_3107 = 9'h82 == T_24222 ? T_48687_130 : GEN_3106;
  assign GEN_3108 = 9'h83 == T_24222 ? T_48687_131 : GEN_3107;
  assign GEN_3109 = 9'h84 == T_24222 ? T_48687_132 : GEN_3108;
  assign GEN_3110 = 9'h85 == T_24222 ? T_48687_133 : GEN_3109;
  assign GEN_3111 = 9'h86 == T_24222 ? T_48687_134 : GEN_3110;
  assign GEN_3112 = 9'h87 == T_24222 ? T_48687_135 : GEN_3111;
  assign GEN_3113 = 9'h88 == T_24222 ? T_48687_136 : GEN_3112;
  assign GEN_3114 = 9'h89 == T_24222 ? T_48687_137 : GEN_3113;
  assign GEN_3115 = 9'h8a == T_24222 ? T_48687_138 : GEN_3114;
  assign GEN_3116 = 9'h8b == T_24222 ? T_48687_139 : GEN_3115;
  assign GEN_3117 = 9'h8c == T_24222 ? T_48687_140 : GEN_3116;
  assign GEN_3118 = 9'h8d == T_24222 ? T_48687_141 : GEN_3117;
  assign GEN_3119 = 9'h8e == T_24222 ? T_48687_142 : GEN_3118;
  assign GEN_3120 = 9'h8f == T_24222 ? T_48687_143 : GEN_3119;
  assign GEN_3121 = 9'h90 == T_24222 ? T_48687_144 : GEN_3120;
  assign GEN_3122 = 9'h91 == T_24222 ? T_48687_145 : GEN_3121;
  assign GEN_3123 = 9'h92 == T_24222 ? T_48687_146 : GEN_3122;
  assign GEN_3124 = 9'h93 == T_24222 ? T_48687_147 : GEN_3123;
  assign GEN_3125 = 9'h94 == T_24222 ? T_48687_148 : GEN_3124;
  assign GEN_3126 = 9'h95 == T_24222 ? T_48687_149 : GEN_3125;
  assign GEN_3127 = 9'h96 == T_24222 ? T_48687_150 : GEN_3126;
  assign GEN_3128 = 9'h97 == T_24222 ? T_48687_151 : GEN_3127;
  assign GEN_3129 = 9'h98 == T_24222 ? T_48687_152 : GEN_3128;
  assign GEN_3130 = 9'h99 == T_24222 ? T_48687_153 : GEN_3129;
  assign GEN_3131 = 9'h9a == T_24222 ? T_48687_154 : GEN_3130;
  assign GEN_3132 = 9'h9b == T_24222 ? T_48687_155 : GEN_3131;
  assign GEN_3133 = 9'h9c == T_24222 ? T_48687_156 : GEN_3132;
  assign GEN_3134 = 9'h9d == T_24222 ? T_48687_157 : GEN_3133;
  assign GEN_3135 = 9'h9e == T_24222 ? T_48687_158 : GEN_3134;
  assign GEN_3136 = 9'h9f == T_24222 ? T_48687_159 : GEN_3135;
  assign GEN_3137 = 9'ha0 == T_24222 ? T_48687_160 : GEN_3136;
  assign GEN_3138 = 9'ha1 == T_24222 ? T_48687_161 : GEN_3137;
  assign GEN_3139 = 9'ha2 == T_24222 ? T_48687_162 : GEN_3138;
  assign GEN_3140 = 9'ha3 == T_24222 ? T_48687_163 : GEN_3139;
  assign GEN_3141 = 9'ha4 == T_24222 ? T_48687_164 : GEN_3140;
  assign GEN_3142 = 9'ha5 == T_24222 ? T_48687_165 : GEN_3141;
  assign GEN_3143 = 9'ha6 == T_24222 ? T_48687_166 : GEN_3142;
  assign GEN_3144 = 9'ha7 == T_24222 ? T_48687_167 : GEN_3143;
  assign GEN_3145 = 9'ha8 == T_24222 ? T_48687_168 : GEN_3144;
  assign GEN_3146 = 9'ha9 == T_24222 ? T_48687_169 : GEN_3145;
  assign GEN_3147 = 9'haa == T_24222 ? T_48687_170 : GEN_3146;
  assign GEN_3148 = 9'hab == T_24222 ? T_48687_171 : GEN_3147;
  assign GEN_3149 = 9'hac == T_24222 ? T_48687_172 : GEN_3148;
  assign GEN_3150 = 9'had == T_24222 ? T_48687_173 : GEN_3149;
  assign GEN_3151 = 9'hae == T_24222 ? T_48687_174 : GEN_3150;
  assign GEN_3152 = 9'haf == T_24222 ? T_48687_175 : GEN_3151;
  assign GEN_3153 = 9'hb0 == T_24222 ? T_48687_176 : GEN_3152;
  assign GEN_3154 = 9'hb1 == T_24222 ? T_48687_177 : GEN_3153;
  assign GEN_3155 = 9'hb2 == T_24222 ? T_48687_178 : GEN_3154;
  assign GEN_3156 = 9'hb3 == T_24222 ? T_48687_179 : GEN_3155;
  assign GEN_3157 = 9'hb4 == T_24222 ? T_48687_180 : GEN_3156;
  assign GEN_3158 = 9'hb5 == T_24222 ? T_48687_181 : GEN_3157;
  assign GEN_3159 = 9'hb6 == T_24222 ? T_48687_182 : GEN_3158;
  assign GEN_3160 = 9'hb7 == T_24222 ? T_48687_183 : GEN_3159;
  assign GEN_3161 = 9'hb8 == T_24222 ? T_48687_184 : GEN_3160;
  assign GEN_3162 = 9'hb9 == T_24222 ? T_48687_185 : GEN_3161;
  assign GEN_3163 = 9'hba == T_24222 ? T_48687_186 : GEN_3162;
  assign GEN_3164 = 9'hbb == T_24222 ? T_48687_187 : GEN_3163;
  assign GEN_3165 = 9'hbc == T_24222 ? T_48687_188 : GEN_3164;
  assign GEN_3166 = 9'hbd == T_24222 ? T_48687_189 : GEN_3165;
  assign GEN_3167 = 9'hbe == T_24222 ? T_48687_190 : GEN_3166;
  assign GEN_3168 = 9'hbf == T_24222 ? T_48687_191 : GEN_3167;
  assign GEN_3169 = 9'hc0 == T_24222 ? T_48687_192 : GEN_3168;
  assign GEN_3170 = 9'hc1 == T_24222 ? T_48687_193 : GEN_3169;
  assign GEN_3171 = 9'hc2 == T_24222 ? T_48687_194 : GEN_3170;
  assign GEN_3172 = 9'hc3 == T_24222 ? T_48687_195 : GEN_3171;
  assign GEN_3173 = 9'hc4 == T_24222 ? T_48687_196 : GEN_3172;
  assign GEN_3174 = 9'hc5 == T_24222 ? T_48687_197 : GEN_3173;
  assign GEN_3175 = 9'hc6 == T_24222 ? T_48687_198 : GEN_3174;
  assign GEN_3176 = 9'hc7 == T_24222 ? T_48687_199 : GEN_3175;
  assign GEN_3177 = 9'hc8 == T_24222 ? T_48687_200 : GEN_3176;
  assign GEN_3178 = 9'hc9 == T_24222 ? T_48687_201 : GEN_3177;
  assign GEN_3179 = 9'hca == T_24222 ? T_48687_202 : GEN_3178;
  assign GEN_3180 = 9'hcb == T_24222 ? T_48687_203 : GEN_3179;
  assign GEN_3181 = 9'hcc == T_24222 ? T_48687_204 : GEN_3180;
  assign GEN_3182 = 9'hcd == T_24222 ? T_48687_205 : GEN_3181;
  assign GEN_3183 = 9'hce == T_24222 ? T_48687_206 : GEN_3182;
  assign GEN_3184 = 9'hcf == T_24222 ? T_48687_207 : GEN_3183;
  assign GEN_3185 = 9'hd0 == T_24222 ? T_48687_208 : GEN_3184;
  assign GEN_3186 = 9'hd1 == T_24222 ? T_48687_209 : GEN_3185;
  assign GEN_3187 = 9'hd2 == T_24222 ? T_48687_210 : GEN_3186;
  assign GEN_3188 = 9'hd3 == T_24222 ? T_48687_211 : GEN_3187;
  assign GEN_3189 = 9'hd4 == T_24222 ? T_48687_212 : GEN_3188;
  assign GEN_3190 = 9'hd5 == T_24222 ? T_48687_213 : GEN_3189;
  assign GEN_3191 = 9'hd6 == T_24222 ? T_48687_214 : GEN_3190;
  assign GEN_3192 = 9'hd7 == T_24222 ? T_48687_215 : GEN_3191;
  assign GEN_3193 = 9'hd8 == T_24222 ? T_48687_216 : GEN_3192;
  assign GEN_3194 = 9'hd9 == T_24222 ? T_48687_217 : GEN_3193;
  assign GEN_3195 = 9'hda == T_24222 ? T_48687_218 : GEN_3194;
  assign GEN_3196 = 9'hdb == T_24222 ? T_48687_219 : GEN_3195;
  assign GEN_3197 = 9'hdc == T_24222 ? T_48687_220 : GEN_3196;
  assign GEN_3198 = 9'hdd == T_24222 ? T_48687_221 : GEN_3197;
  assign GEN_3199 = 9'hde == T_24222 ? T_48687_222 : GEN_3198;
  assign GEN_3200 = 9'hdf == T_24222 ? T_48687_223 : GEN_3199;
  assign GEN_3201 = 9'he0 == T_24222 ? T_48687_224 : GEN_3200;
  assign GEN_3202 = 9'he1 == T_24222 ? T_48687_225 : GEN_3201;
  assign GEN_3203 = 9'he2 == T_24222 ? T_48687_226 : GEN_3202;
  assign GEN_3204 = 9'he3 == T_24222 ? T_48687_227 : GEN_3203;
  assign GEN_3205 = 9'he4 == T_24222 ? T_48687_228 : GEN_3204;
  assign GEN_3206 = 9'he5 == T_24222 ? T_48687_229 : GEN_3205;
  assign GEN_3207 = 9'he6 == T_24222 ? T_48687_230 : GEN_3206;
  assign GEN_3208 = 9'he7 == T_24222 ? T_48687_231 : GEN_3207;
  assign GEN_3209 = 9'he8 == T_24222 ? T_48687_232 : GEN_3208;
  assign GEN_3210 = 9'he9 == T_24222 ? T_48687_233 : GEN_3209;
  assign GEN_3211 = 9'hea == T_24222 ? T_48687_234 : GEN_3210;
  assign GEN_3212 = 9'heb == T_24222 ? T_48687_235 : GEN_3211;
  assign GEN_3213 = 9'hec == T_24222 ? T_48687_236 : GEN_3212;
  assign GEN_3214 = 9'hed == T_24222 ? T_48687_237 : GEN_3213;
  assign GEN_3215 = 9'hee == T_24222 ? T_48687_238 : GEN_3214;
  assign GEN_3216 = 9'hef == T_24222 ? T_48687_239 : GEN_3215;
  assign GEN_3217 = 9'hf0 == T_24222 ? T_48687_240 : GEN_3216;
  assign GEN_3218 = 9'hf1 == T_24222 ? T_48687_241 : GEN_3217;
  assign GEN_3219 = 9'hf2 == T_24222 ? T_48687_242 : GEN_3218;
  assign GEN_3220 = 9'hf3 == T_24222 ? T_48687_243 : GEN_3219;
  assign GEN_3221 = 9'hf4 == T_24222 ? T_48687_244 : GEN_3220;
  assign GEN_3222 = 9'hf5 == T_24222 ? T_48687_245 : GEN_3221;
  assign GEN_3223 = 9'hf6 == T_24222 ? T_48687_246 : GEN_3222;
  assign GEN_3224 = 9'hf7 == T_24222 ? T_48687_247 : GEN_3223;
  assign GEN_3225 = 9'hf8 == T_24222 ? T_48687_248 : GEN_3224;
  assign GEN_3226 = 9'hf9 == T_24222 ? T_48687_249 : GEN_3225;
  assign GEN_3227 = 9'hfa == T_24222 ? T_48687_250 : GEN_3226;
  assign GEN_3228 = 9'hfb == T_24222 ? T_48687_251 : GEN_3227;
  assign GEN_3229 = 9'hfc == T_24222 ? T_48687_252 : GEN_3228;
  assign GEN_3230 = 9'hfd == T_24222 ? T_48687_253 : GEN_3229;
  assign GEN_3231 = 9'hfe == T_24222 ? T_48687_254 : GEN_3230;
  assign GEN_3232 = 9'hff == T_24222 ? T_48687_255 : GEN_3231;
  assign GEN_3233 = 9'h100 == T_24222 ? T_48687_256 : GEN_3232;
  assign GEN_3234 = 9'h101 == T_24222 ? T_48687_257 : GEN_3233;
  assign GEN_3235 = 9'h102 == T_24222 ? T_48687_258 : GEN_3234;
  assign GEN_3236 = 9'h103 == T_24222 ? T_48687_259 : GEN_3235;
  assign GEN_3237 = 9'h104 == T_24222 ? T_48687_260 : GEN_3236;
  assign GEN_3238 = 9'h105 == T_24222 ? T_48687_261 : GEN_3237;
  assign GEN_3239 = 9'h106 == T_24222 ? T_48687_262 : GEN_3238;
  assign GEN_3240 = 9'h107 == T_24222 ? T_48687_263 : GEN_3239;
  assign GEN_3241 = 9'h108 == T_24222 ? T_48687_264 : GEN_3240;
  assign GEN_3242 = 9'h109 == T_24222 ? T_48687_265 : GEN_3241;
  assign GEN_3243 = 9'h10a == T_24222 ? T_48687_266 : GEN_3242;
  assign GEN_3244 = 9'h10b == T_24222 ? T_48687_267 : GEN_3243;
  assign GEN_3245 = 9'h10c == T_24222 ? T_48687_268 : GEN_3244;
  assign GEN_3246 = 9'h10d == T_24222 ? T_48687_269 : GEN_3245;
  assign GEN_3247 = 9'h10e == T_24222 ? T_48687_270 : GEN_3246;
  assign GEN_3248 = 9'h10f == T_24222 ? T_48687_271 : GEN_3247;
  assign GEN_3249 = 9'h110 == T_24222 ? T_48687_272 : GEN_3248;
  assign GEN_3250 = 9'h111 == T_24222 ? T_48687_273 : GEN_3249;
  assign GEN_3251 = 9'h112 == T_24222 ? T_48687_274 : GEN_3250;
  assign GEN_3252 = 9'h113 == T_24222 ? T_48687_275 : GEN_3251;
  assign GEN_3253 = 9'h114 == T_24222 ? T_48687_276 : GEN_3252;
  assign GEN_3254 = 9'h115 == T_24222 ? T_48687_277 : GEN_3253;
  assign GEN_3255 = 9'h116 == T_24222 ? T_48687_278 : GEN_3254;
  assign GEN_3256 = 9'h117 == T_24222 ? T_48687_279 : GEN_3255;
  assign GEN_3257 = 9'h118 == T_24222 ? T_48687_280 : GEN_3256;
  assign GEN_3258 = 9'h119 == T_24222 ? T_48687_281 : GEN_3257;
  assign GEN_3259 = 9'h11a == T_24222 ? T_48687_282 : GEN_3258;
  assign GEN_3260 = 9'h11b == T_24222 ? T_48687_283 : GEN_3259;
  assign GEN_3261 = 9'h11c == T_24222 ? T_48687_284 : GEN_3260;
  assign GEN_3262 = 9'h11d == T_24222 ? T_48687_285 : GEN_3261;
  assign GEN_3263 = 9'h11e == T_24222 ? T_48687_286 : GEN_3262;
  assign GEN_3264 = 9'h11f == T_24222 ? T_48687_287 : GEN_3263;
  assign GEN_3265 = 9'h120 == T_24222 ? T_48687_288 : GEN_3264;
  assign GEN_3266 = 9'h121 == T_24222 ? T_48687_289 : GEN_3265;
  assign GEN_3267 = 9'h122 == T_24222 ? T_48687_290 : GEN_3266;
  assign GEN_3268 = 9'h123 == T_24222 ? T_48687_291 : GEN_3267;
  assign GEN_3269 = 9'h124 == T_24222 ? T_48687_292 : GEN_3268;
  assign GEN_3270 = 9'h125 == T_24222 ? T_48687_293 : GEN_3269;
  assign GEN_3271 = 9'h126 == T_24222 ? T_48687_294 : GEN_3270;
  assign GEN_3272 = 9'h127 == T_24222 ? T_48687_295 : GEN_3271;
  assign GEN_3273 = 9'h128 == T_24222 ? T_48687_296 : GEN_3272;
  assign GEN_3274 = 9'h129 == T_24222 ? T_48687_297 : GEN_3273;
  assign GEN_3275 = 9'h12a == T_24222 ? T_48687_298 : GEN_3274;
  assign GEN_3276 = 9'h12b == T_24222 ? T_48687_299 : GEN_3275;
  assign GEN_3277 = 9'h12c == T_24222 ? T_48687_300 : GEN_3276;
  assign GEN_3278 = 9'h12d == T_24222 ? T_48687_301 : GEN_3277;
  assign GEN_3279 = 9'h12e == T_24222 ? T_48687_302 : GEN_3278;
  assign GEN_3280 = 9'h12f == T_24222 ? T_48687_303 : GEN_3279;
  assign GEN_3281 = 9'h130 == T_24222 ? T_48687_304 : GEN_3280;
  assign GEN_3282 = 9'h131 == T_24222 ? T_48687_305 : GEN_3281;
  assign GEN_3283 = 9'h132 == T_24222 ? T_48687_306 : GEN_3282;
  assign GEN_3284 = 9'h133 == T_24222 ? T_48687_307 : GEN_3283;
  assign GEN_3285 = 9'h134 == T_24222 ? T_48687_308 : GEN_3284;
  assign GEN_3286 = 9'h135 == T_24222 ? T_48687_309 : GEN_3285;
  assign GEN_3287 = 9'h136 == T_24222 ? T_48687_310 : GEN_3286;
  assign GEN_3288 = 9'h137 == T_24222 ? T_48687_311 : GEN_3287;
  assign GEN_3289 = 9'h138 == T_24222 ? T_48687_312 : GEN_3288;
  assign GEN_3290 = 9'h139 == T_24222 ? T_48687_313 : GEN_3289;
  assign GEN_3291 = 9'h13a == T_24222 ? T_48687_314 : GEN_3290;
  assign GEN_3292 = 9'h13b == T_24222 ? T_48687_315 : GEN_3291;
  assign GEN_3293 = 9'h13c == T_24222 ? T_48687_316 : GEN_3292;
  assign GEN_3294 = 9'h13d == T_24222 ? T_48687_317 : GEN_3293;
  assign GEN_3295 = 9'h13e == T_24222 ? T_48687_318 : GEN_3294;
  assign GEN_3296 = 9'h13f == T_24222 ? T_48687_319 : GEN_3295;
  assign GEN_3297 = 9'h140 == T_24222 ? T_48687_320 : GEN_3296;
  assign GEN_3298 = 9'h141 == T_24222 ? T_48687_321 : GEN_3297;
  assign GEN_3299 = 9'h142 == T_24222 ? T_48687_322 : GEN_3298;
  assign GEN_3300 = 9'h143 == T_24222 ? T_48687_323 : GEN_3299;
  assign GEN_3301 = 9'h144 == T_24222 ? T_48687_324 : GEN_3300;
  assign GEN_3302 = 9'h145 == T_24222 ? T_48687_325 : GEN_3301;
  assign GEN_3303 = 9'h146 == T_24222 ? T_48687_326 : GEN_3302;
  assign GEN_3304 = 9'h147 == T_24222 ? T_48687_327 : GEN_3303;
  assign GEN_3305 = 9'h148 == T_24222 ? T_48687_328 : GEN_3304;
  assign GEN_3306 = 9'h149 == T_24222 ? T_48687_329 : GEN_3305;
  assign GEN_3307 = 9'h14a == T_24222 ? T_48687_330 : GEN_3306;
  assign GEN_3308 = 9'h14b == T_24222 ? T_48687_331 : GEN_3307;
  assign GEN_3309 = 9'h14c == T_24222 ? T_48687_332 : GEN_3308;
  assign GEN_3310 = 9'h14d == T_24222 ? T_48687_333 : GEN_3309;
  assign GEN_3311 = 9'h14e == T_24222 ? T_48687_334 : GEN_3310;
  assign GEN_3312 = 9'h14f == T_24222 ? T_48687_335 : GEN_3311;
  assign GEN_3313 = 9'h150 == T_24222 ? T_48687_336 : GEN_3312;
  assign GEN_3314 = 9'h151 == T_24222 ? T_48687_337 : GEN_3313;
  assign GEN_3315 = 9'h152 == T_24222 ? T_48687_338 : GEN_3314;
  assign GEN_3316 = 9'h153 == T_24222 ? T_48687_339 : GEN_3315;
  assign GEN_3317 = 9'h154 == T_24222 ? T_48687_340 : GEN_3316;
  assign GEN_3318 = 9'h155 == T_24222 ? T_48687_341 : GEN_3317;
  assign GEN_3319 = 9'h156 == T_24222 ? T_48687_342 : GEN_3318;
  assign GEN_3320 = 9'h157 == T_24222 ? T_48687_343 : GEN_3319;
  assign GEN_3321 = 9'h158 == T_24222 ? T_48687_344 : GEN_3320;
  assign GEN_3322 = 9'h159 == T_24222 ? T_48687_345 : GEN_3321;
  assign GEN_3323 = 9'h15a == T_24222 ? T_48687_346 : GEN_3322;
  assign GEN_3324 = 9'h15b == T_24222 ? T_48687_347 : GEN_3323;
  assign GEN_3325 = 9'h15c == T_24222 ? T_48687_348 : GEN_3324;
  assign GEN_3326 = 9'h15d == T_24222 ? T_48687_349 : GEN_3325;
  assign GEN_3327 = 9'h15e == T_24222 ? T_48687_350 : GEN_3326;
  assign GEN_3328 = 9'h15f == T_24222 ? T_48687_351 : GEN_3327;
  assign GEN_3329 = 9'h160 == T_24222 ? T_48687_352 : GEN_3328;
  assign GEN_3330 = 9'h161 == T_24222 ? T_48687_353 : GEN_3329;
  assign GEN_3331 = 9'h162 == T_24222 ? T_48687_354 : GEN_3330;
  assign GEN_3332 = 9'h163 == T_24222 ? T_48687_355 : GEN_3331;
  assign GEN_3333 = 9'h164 == T_24222 ? T_48687_356 : GEN_3332;
  assign GEN_3334 = 9'h165 == T_24222 ? T_48687_357 : GEN_3333;
  assign GEN_3335 = 9'h166 == T_24222 ? T_48687_358 : GEN_3334;
  assign GEN_3336 = 9'h167 == T_24222 ? T_48687_359 : GEN_3335;
  assign GEN_3337 = 9'h168 == T_24222 ? T_48687_360 : GEN_3336;
  assign GEN_3338 = 9'h169 == T_24222 ? T_48687_361 : GEN_3337;
  assign GEN_3339 = 9'h16a == T_24222 ? T_48687_362 : GEN_3338;
  assign GEN_3340 = 9'h16b == T_24222 ? T_48687_363 : GEN_3339;
  assign GEN_3341 = 9'h16c == T_24222 ? T_48687_364 : GEN_3340;
  assign GEN_3342 = 9'h16d == T_24222 ? T_48687_365 : GEN_3341;
  assign GEN_3343 = 9'h16e == T_24222 ? T_48687_366 : GEN_3342;
  assign GEN_3344 = 9'h16f == T_24222 ? T_48687_367 : GEN_3343;
  assign GEN_3345 = 9'h170 == T_24222 ? T_48687_368 : GEN_3344;
  assign GEN_3346 = 9'h171 == T_24222 ? T_48687_369 : GEN_3345;
  assign GEN_3347 = 9'h172 == T_24222 ? T_48687_370 : GEN_3346;
  assign GEN_3348 = 9'h173 == T_24222 ? T_48687_371 : GEN_3347;
  assign GEN_3349 = 9'h174 == T_24222 ? T_48687_372 : GEN_3348;
  assign GEN_3350 = 9'h175 == T_24222 ? T_48687_373 : GEN_3349;
  assign GEN_3351 = 9'h176 == T_24222 ? T_48687_374 : GEN_3350;
  assign GEN_3352 = 9'h177 == T_24222 ? T_48687_375 : GEN_3351;
  assign GEN_3353 = 9'h178 == T_24222 ? T_48687_376 : GEN_3352;
  assign GEN_3354 = 9'h179 == T_24222 ? T_48687_377 : GEN_3353;
  assign GEN_3355 = 9'h17a == T_24222 ? T_48687_378 : GEN_3354;
  assign GEN_3356 = 9'h17b == T_24222 ? T_48687_379 : GEN_3355;
  assign GEN_3357 = 9'h17c == T_24222 ? T_48687_380 : GEN_3356;
  assign GEN_3358 = 9'h17d == T_24222 ? T_48687_381 : GEN_3357;
  assign GEN_3359 = 9'h17e == T_24222 ? T_48687_382 : GEN_3358;
  assign GEN_3360 = 9'h17f == T_24222 ? T_48687_383 : GEN_3359;
  assign GEN_3361 = 9'h180 == T_24222 ? T_48687_384 : GEN_3360;
  assign GEN_3362 = 9'h181 == T_24222 ? T_48687_385 : GEN_3361;
  assign GEN_3363 = 9'h182 == T_24222 ? T_48687_386 : GEN_3362;
  assign GEN_3364 = 9'h183 == T_24222 ? T_48687_387 : GEN_3363;
  assign GEN_3365 = 9'h184 == T_24222 ? T_48687_388 : GEN_3364;
  assign GEN_3366 = 9'h185 == T_24222 ? T_48687_389 : GEN_3365;
  assign GEN_3367 = 9'h186 == T_24222 ? T_48687_390 : GEN_3366;
  assign GEN_3368 = 9'h187 == T_24222 ? T_48687_391 : GEN_3367;
  assign GEN_3369 = 9'h188 == T_24222 ? T_48687_392 : GEN_3368;
  assign GEN_3370 = 9'h189 == T_24222 ? T_48687_393 : GEN_3369;
  assign GEN_3371 = 9'h18a == T_24222 ? T_48687_394 : GEN_3370;
  assign GEN_3372 = 9'h18b == T_24222 ? T_48687_395 : GEN_3371;
  assign GEN_3373 = 9'h18c == T_24222 ? T_48687_396 : GEN_3372;
  assign GEN_3374 = 9'h18d == T_24222 ? T_48687_397 : GEN_3373;
  assign GEN_3375 = 9'h18e == T_24222 ? T_48687_398 : GEN_3374;
  assign GEN_3376 = 9'h18f == T_24222 ? T_48687_399 : GEN_3375;
  assign GEN_3377 = 9'h190 == T_24222 ? T_48687_400 : GEN_3376;
  assign GEN_3378 = 9'h191 == T_24222 ? T_48687_401 : GEN_3377;
  assign GEN_3379 = 9'h192 == T_24222 ? T_48687_402 : GEN_3378;
  assign GEN_3380 = 9'h193 == T_24222 ? T_48687_403 : GEN_3379;
  assign GEN_3381 = 9'h194 == T_24222 ? T_48687_404 : GEN_3380;
  assign GEN_3382 = 9'h195 == T_24222 ? T_48687_405 : GEN_3381;
  assign GEN_3383 = 9'h196 == T_24222 ? T_48687_406 : GEN_3382;
  assign GEN_3384 = 9'h197 == T_24222 ? T_48687_407 : GEN_3383;
  assign GEN_3385 = 9'h198 == T_24222 ? T_48687_408 : GEN_3384;
  assign GEN_3386 = 9'h199 == T_24222 ? T_48687_409 : GEN_3385;
  assign GEN_3387 = 9'h19a == T_24222 ? T_48687_410 : GEN_3386;
  assign GEN_3388 = 9'h19b == T_24222 ? T_48687_411 : GEN_3387;
  assign GEN_3389 = 9'h19c == T_24222 ? T_48687_412 : GEN_3388;
  assign GEN_3390 = 9'h19d == T_24222 ? T_48687_413 : GEN_3389;
  assign GEN_3391 = 9'h19e == T_24222 ? T_48687_414 : GEN_3390;
  assign GEN_3392 = 9'h19f == T_24222 ? T_48687_415 : GEN_3391;
  assign GEN_3393 = 9'h1a0 == T_24222 ? T_48687_416 : GEN_3392;
  assign GEN_3394 = 9'h1a1 == T_24222 ? T_48687_417 : GEN_3393;
  assign GEN_3395 = 9'h1a2 == T_24222 ? T_48687_418 : GEN_3394;
  assign GEN_3396 = 9'h1a3 == T_24222 ? T_48687_419 : GEN_3395;
  assign GEN_3397 = 9'h1a4 == T_24222 ? T_48687_420 : GEN_3396;
  assign GEN_3398 = 9'h1a5 == T_24222 ? T_48687_421 : GEN_3397;
  assign GEN_3399 = 9'h1a6 == T_24222 ? T_48687_422 : GEN_3398;
  assign GEN_3400 = 9'h1a7 == T_24222 ? T_48687_423 : GEN_3399;
  assign GEN_3401 = 9'h1a8 == T_24222 ? T_48687_424 : GEN_3400;
  assign GEN_3402 = 9'h1a9 == T_24222 ? T_48687_425 : GEN_3401;
  assign GEN_3403 = 9'h1aa == T_24222 ? T_48687_426 : GEN_3402;
  assign GEN_3404 = 9'h1ab == T_24222 ? T_48687_427 : GEN_3403;
  assign GEN_3405 = 9'h1ac == T_24222 ? T_48687_428 : GEN_3404;
  assign GEN_3406 = 9'h1ad == T_24222 ? T_48687_429 : GEN_3405;
  assign GEN_3407 = 9'h1ae == T_24222 ? T_48687_430 : GEN_3406;
  assign GEN_3408 = 9'h1af == T_24222 ? T_48687_431 : GEN_3407;
  assign GEN_3409 = 9'h1b0 == T_24222 ? T_48687_432 : GEN_3408;
  assign GEN_3410 = 9'h1b1 == T_24222 ? T_48687_433 : GEN_3409;
  assign GEN_3411 = 9'h1b2 == T_24222 ? T_48687_434 : GEN_3410;
  assign GEN_3412 = 9'h1b3 == T_24222 ? T_48687_435 : GEN_3411;
  assign GEN_3413 = 9'h1b4 == T_24222 ? T_48687_436 : GEN_3412;
  assign GEN_3414 = 9'h1b5 == T_24222 ? T_48687_437 : GEN_3413;
  assign GEN_3415 = 9'h1b6 == T_24222 ? T_48687_438 : GEN_3414;
  assign GEN_3416 = 9'h1b7 == T_24222 ? T_48687_439 : GEN_3415;
  assign GEN_3417 = 9'h1b8 == T_24222 ? T_48687_440 : GEN_3416;
  assign GEN_3418 = 9'h1b9 == T_24222 ? T_48687_441 : GEN_3417;
  assign GEN_3419 = 9'h1ba == T_24222 ? T_48687_442 : GEN_3418;
  assign GEN_3420 = 9'h1bb == T_24222 ? T_48687_443 : GEN_3419;
  assign GEN_3421 = 9'h1bc == T_24222 ? T_48687_444 : GEN_3420;
  assign GEN_3422 = 9'h1bd == T_24222 ? T_48687_445 : GEN_3421;
  assign GEN_3423 = 9'h1be == T_24222 ? T_48687_446 : GEN_3422;
  assign GEN_3424 = 9'h1bf == T_24222 ? T_48687_447 : GEN_3423;
  assign GEN_3425 = 9'h1c0 == T_24222 ? T_48687_448 : GEN_3424;
  assign GEN_3426 = 9'h1c1 == T_24222 ? T_48687_449 : GEN_3425;
  assign GEN_3427 = 9'h1c2 == T_24222 ? T_48687_450 : GEN_3426;
  assign GEN_3428 = 9'h1c3 == T_24222 ? T_48687_451 : GEN_3427;
  assign GEN_3429 = 9'h1c4 == T_24222 ? T_48687_452 : GEN_3428;
  assign GEN_3430 = 9'h1c5 == T_24222 ? T_48687_453 : GEN_3429;
  assign GEN_3431 = 9'h1c6 == T_24222 ? T_48687_454 : GEN_3430;
  assign GEN_3432 = 9'h1c7 == T_24222 ? T_48687_455 : GEN_3431;
  assign GEN_3433 = 9'h1c8 == T_24222 ? T_48687_456 : GEN_3432;
  assign GEN_3434 = 9'h1c9 == T_24222 ? T_48687_457 : GEN_3433;
  assign GEN_3435 = 9'h1ca == T_24222 ? T_48687_458 : GEN_3434;
  assign GEN_3436 = 9'h1cb == T_24222 ? T_48687_459 : GEN_3435;
  assign GEN_3437 = 9'h1cc == T_24222 ? T_48687_460 : GEN_3436;
  assign GEN_3438 = 9'h1cd == T_24222 ? T_48687_461 : GEN_3437;
  assign GEN_3439 = 9'h1ce == T_24222 ? T_48687_462 : GEN_3438;
  assign GEN_3440 = 9'h1cf == T_24222 ? T_48687_463 : GEN_3439;
  assign GEN_3441 = 9'h1d0 == T_24222 ? T_48687_464 : GEN_3440;
  assign GEN_3442 = 9'h1d1 == T_24222 ? T_48687_465 : GEN_3441;
  assign GEN_3443 = 9'h1d2 == T_24222 ? T_48687_466 : GEN_3442;
  assign GEN_3444 = 9'h1d3 == T_24222 ? T_48687_467 : GEN_3443;
  assign GEN_3445 = 9'h1d4 == T_24222 ? T_48687_468 : GEN_3444;
  assign GEN_3446 = 9'h1d5 == T_24222 ? T_48687_469 : GEN_3445;
  assign GEN_3447 = 9'h1d6 == T_24222 ? T_48687_470 : GEN_3446;
  assign GEN_3448 = 9'h1d7 == T_24222 ? T_48687_471 : GEN_3447;
  assign GEN_3449 = 9'h1d8 == T_24222 ? T_48687_472 : GEN_3448;
  assign GEN_3450 = 9'h1d9 == T_24222 ? T_48687_473 : GEN_3449;
  assign GEN_3451 = 9'h1da == T_24222 ? T_48687_474 : GEN_3450;
  assign GEN_3452 = 9'h1db == T_24222 ? T_48687_475 : GEN_3451;
  assign GEN_3453 = 9'h1dc == T_24222 ? T_48687_476 : GEN_3452;
  assign GEN_3454 = 9'h1dd == T_24222 ? T_48687_477 : GEN_3453;
  assign GEN_3455 = 9'h1de == T_24222 ? T_48687_478 : GEN_3454;
  assign GEN_3456 = 9'h1df == T_24222 ? T_48687_479 : GEN_3455;
  assign GEN_3457 = 9'h1e0 == T_24222 ? T_48687_480 : GEN_3456;
  assign GEN_3458 = 9'h1e1 == T_24222 ? T_48687_481 : GEN_3457;
  assign GEN_3459 = 9'h1e2 == T_24222 ? T_48687_482 : GEN_3458;
  assign GEN_3460 = 9'h1e3 == T_24222 ? T_48687_483 : GEN_3459;
  assign GEN_3461 = 9'h1e4 == T_24222 ? T_48687_484 : GEN_3460;
  assign GEN_3462 = 9'h1e5 == T_24222 ? T_48687_485 : GEN_3461;
  assign GEN_3463 = 9'h1e6 == T_24222 ? T_48687_486 : GEN_3462;
  assign GEN_3464 = 9'h1e7 == T_24222 ? T_48687_487 : GEN_3463;
  assign GEN_3465 = 9'h1e8 == T_24222 ? T_48687_488 : GEN_3464;
  assign GEN_3466 = 9'h1e9 == T_24222 ? T_48687_489 : GEN_3465;
  assign GEN_3467 = 9'h1ea == T_24222 ? T_48687_490 : GEN_3466;
  assign GEN_3468 = 9'h1eb == T_24222 ? T_48687_491 : GEN_3467;
  assign GEN_3469 = 9'h1ec == T_24222 ? T_48687_492 : GEN_3468;
  assign GEN_3470 = 9'h1ed == T_24222 ? T_48687_493 : GEN_3469;
  assign GEN_3471 = 9'h1ee == T_24222 ? T_48687_494 : GEN_3470;
  assign GEN_3472 = 9'h1ef == T_24222 ? T_48687_495 : GEN_3471;
  assign GEN_3473 = 9'h1f0 == T_24222 ? T_48687_496 : GEN_3472;
  assign GEN_3474 = 9'h1f1 == T_24222 ? T_48687_497 : GEN_3473;
  assign GEN_3475 = 9'h1f2 == T_24222 ? T_48687_498 : GEN_3474;
  assign GEN_3476 = 9'h1f3 == T_24222 ? T_48687_499 : GEN_3475;
  assign GEN_3477 = 9'h1f4 == T_24222 ? T_48687_500 : GEN_3476;
  assign GEN_3478 = 9'h1f5 == T_24222 ? T_48687_501 : GEN_3477;
  assign GEN_3479 = 9'h1f6 == T_24222 ? T_48687_502 : GEN_3478;
  assign GEN_3480 = 9'h1f7 == T_24222 ? T_48687_503 : GEN_3479;
  assign GEN_3481 = 9'h1f8 == T_24222 ? T_48687_504 : GEN_3480;
  assign GEN_3482 = 9'h1f9 == T_24222 ? T_48687_505 : GEN_3481;
  assign GEN_3483 = 9'h1fa == T_24222 ? T_48687_506 : GEN_3482;
  assign GEN_3484 = 9'h1fb == T_24222 ? T_48687_507 : GEN_3483;
  assign GEN_3485 = 9'h1fc == T_24222 ? T_48687_508 : GEN_3484;
  assign GEN_3486 = 9'h1fd == T_24222 ? T_48687_509 : GEN_3485;
  assign GEN_3487 = 9'h1fe == T_24222 ? T_48687_510 : GEN_3486;
  assign GEN_3488 = 9'h1ff == T_24222 ? T_48687_511 : GEN_3487;
  assign T_49204 = GEN_7 ? GEN_8 : 32'h0;
  assign T_49205 = T_3169_bits_extra[9:8];
  assign T_49207 = T_3169_bits_extra[7:3];
  assign T_49208 = T_3169_bits_extra[2:0];
  assign T_49219_opcode = 3'h0;
  assign T_49219_param = 2'h0;
  assign T_49219_size = T_49208;
  assign T_49219_source = T_49207;
  assign T_49219_sink = 1'h0;
  assign T_49219_addr_lo = T_49205;
  assign T_49219_data = 32'h0;
  assign T_49219_error = 1'h0;

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      priority_0 <= 3'h0;
      priority_1 <= 3'h0;
      priority_2 <= 3'h0;
      priority_3 <= 3'h0;
      priority_4 <= 3'h0;
      priority_5 <= 3'h0;
      priority_6 <= 3'h0;
      priority_7 <= 3'h0;
      priority_8 <= 3'h0;
      priority_9 <= 3'h0;
      priority_10 <= 3'h0;
      priority_11 <= 3'h0;
      priority_12 <= 3'h0;
      priority_13 <= 3'h0;
      priority_14 <= 3'h0;
      priority_15 <= 3'h0;
      priority_16 <= 3'h0;
      priority_17 <= 3'h0;
      priority_18 <= 3'h0;
      priority_19 <= 3'h0;
      priority_20 <= 3'h0;
      priority_21 <= 3'h0;
      priority_22 <= 3'h0;
      priority_23 <= 3'h0;
      priority_24 <= 3'h0;
      priority_25 <= 3'h0;
      priority_26 <= 3'h0;
      priority_27 <= 3'h0;
      priority_28 <= 3'h0;
      priority_29 <= 3'h0;
      priority_30 <= 3'h0;
      priority_31 <= 3'h0;
      priority_32 <= 3'h0;
      priority_33 <= 3'h0;
      priority_34 <= 3'h0;
      priority_35 <= 3'h0;
      priority_36 <= 3'h0;
      priority_37 <= 3'h0;
      priority_38 <= 3'h0;
      priority_39 <= 3'h0;
      priority_40 <= 3'h0;
      priority_41 <= 3'h0;
      priority_42 <= 3'h0;
      priority_43 <= 3'h0;
      priority_44 <= 3'h0;
      priority_45 <= 3'h0;
      priority_46 <= 3'h0;
      priority_47 <= 3'h0;
      priority_48 <= 3'h0;
      priority_49 <= 3'h0;
      priority_50 <= 3'h0;
      priority_51 <= 3'h0;
      threshold_0 <= 3'h0;
    end
    else begin
      priority_0 <= 3'h0;
      priority_1 <= GEN_349[2:0];
      priority_2 <= GEN_358[2:0];
      priority_3 <= GEN_403[2:0];
      priority_4 <= GEN_420[2:0];
      priority_5 <= GEN_61[2:0];
      priority_6 <= GEN_350[2:0];
      priority_7 <= GEN_401[2:0];
      priority_8 <= GEN_415[2:0];
      priority_9 <= GEN_355[2:0];
      priority_10 <= GEN_62[2:0];
      priority_11 <= GEN_410[2:0];
      priority_12 <= GEN_399[2:0];
      priority_13 <= GEN_356[2:0];
      priority_14 <= GEN_67[2:0];
      priority_15 <= GEN_422[2:0];
      priority_16 <= GEN_408[2:0];
      priority_17 <= GEN_362[2:0];
      priority_18 <= GEN_406[2:0];
      priority_19 <= GEN_419[2:0];
      priority_20 <= GEN_68[2:0];
      priority_21 <= GEN_353[2:0];
      priority_22 <= GEN_396[2:0];
      priority_23 <= GEN_414[2:0];
      priority_24 <= GEN_64[2:0];
      priority_25 <= GEN_66[2:0];
      priority_26 <= GEN_413[2:0];
      priority_27 <= GEN_398[2:0];
      priority_28 <= GEN_351[2:0];
      priority_29 <= GEN_90[2:0];
      priority_30 <= GEN_417[2:0];
      priority_31 <= GEN_409[2:0];
      priority_32 <= GEN_359[2:0];
      priority_33 <= GEN_354[2:0];
      priority_34 <= GEN_360[2:0];
      priority_35 <= GEN_404[2:0];
      priority_36 <= GEN_416[2:0];
      priority_37 <= GEN_65[2:0];
      priority_38 <= GEN_352[2:0];
      priority_39 <= GEN_402[2:0];
      priority_40 <= GEN_412[2:0];
      priority_41 <= GEN_357[2:0];
      priority_42 <= GEN_63[2:0];
      priority_43 <= GEN_411[2:0];
      priority_44 <= GEN_397[2:0];
      priority_45 <= GEN_361[2:0];
      priority_46 <= GEN_89[2:0];
      priority_47 <= GEN_421[2:0];
      priority_48 <= GEN_405[2:0];
      priority_49 <= GEN_400[2:0];
      priority_50 <= GEN_407[2:0];
      priority_51 <= GEN_418[2:0];
      threshold_0 <= GEN_363[2:0];
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_0 <= T_2365_0;
    end else begin
      pending_0 <= 1'h0;
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_1 <= T_2365_1;
    end else begin
      if (T_9487) begin
        if (6'h1 == maxDevs_0) begin
          pending_1 <= GEN_0;
        end else begin
          if (gateways_0_valid) begin
            pending_1 <= 1'h1;
          end
        end
      end else begin
        if (gateways_0_valid) begin
          pending_1 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_2 <= T_2365_2;
    end else begin
      if (T_9487) begin
        if (6'h2 == maxDevs_0) begin
          pending_2 <= GEN_0;
        end else begin
          if (gateways_1_valid) begin
            pending_2 <= 1'h1;
          end
        end
      end else begin
        if (gateways_1_valid) begin
          pending_2 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_3 <= T_2365_3;
    end else begin
      if (T_9487) begin
        if (6'h3 == maxDevs_0) begin
          pending_3 <= GEN_0;
        end else begin
          if (gateways_2_valid) begin
            pending_3 <= 1'h1;
          end
        end
      end else begin
        if (gateways_2_valid) begin
          pending_3 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_4 <= T_2365_4;
    end else begin
      if (T_9487) begin
        if (6'h4 == maxDevs_0) begin
          pending_4 <= GEN_0;
        end else begin
          if (gateways_3_valid) begin
            pending_4 <= 1'h1;
          end
        end
      end else begin
        if (gateways_3_valid) begin
          pending_4 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_5 <= T_2365_5;
    end else begin
      if (T_9487) begin
        if (6'h5 == maxDevs_0) begin
          pending_5 <= GEN_0;
        end else begin
          if (gateways_4_valid) begin
            pending_5 <= 1'h1;
          end
        end
      end else begin
        if (gateways_4_valid) begin
          pending_5 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_6 <= T_2365_6;
    end else begin
      if (T_9487) begin
        if (6'h6 == maxDevs_0) begin
          pending_6 <= GEN_0;
        end else begin
          if (gateways_5_valid) begin
            pending_6 <= 1'h1;
          end
        end
      end else begin
        if (gateways_5_valid) begin
          pending_6 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_7 <= T_2365_7;
    end else begin
      if (T_9487) begin
        if (6'h7 == maxDevs_0) begin
          pending_7 <= GEN_0;
        end else begin
          if (gateways_6_valid) begin
            pending_7 <= 1'h1;
          end
        end
      end else begin
        if (gateways_6_valid) begin
          pending_7 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_8 <= T_2365_8;
    end else begin
      if (T_9487) begin
        if (6'h8 == maxDevs_0) begin
          pending_8 <= GEN_0;
        end else begin
          if (gateways_7_valid) begin
            pending_8 <= 1'h1;
          end
        end
      end else begin
        if (gateways_7_valid) begin
          pending_8 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_9 <= T_2365_9;
    end else begin
      if (T_9487) begin
        if (6'h9 == maxDevs_0) begin
          pending_9 <= GEN_0;
        end else begin
          if (gateways_8_valid) begin
            pending_9 <= 1'h1;
          end
        end
      end else begin
        if (gateways_8_valid) begin
          pending_9 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_10 <= T_2365_10;
    end else begin
      if (T_9487) begin
        if (6'ha == maxDevs_0) begin
          pending_10 <= GEN_0;
        end else begin
          if (gateways_9_valid) begin
            pending_10 <= 1'h1;
          end
        end
      end else begin
        if (gateways_9_valid) begin
          pending_10 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_11 <= T_2365_11;
    end else begin
      if (T_9487) begin
        if (6'hb == maxDevs_0) begin
          pending_11 <= GEN_0;
        end else begin
          if (gateways_10_valid) begin
            pending_11 <= 1'h1;
          end
        end
      end else begin
        if (gateways_10_valid) begin
          pending_11 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_12 <= T_2365_12;
    end else begin
      if (T_9487) begin
        if (6'hc == maxDevs_0) begin
          pending_12 <= GEN_0;
        end else begin
          if (gateways_11_valid) begin
            pending_12 <= 1'h1;
          end
        end
      end else begin
        if (gateways_11_valid) begin
          pending_12 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_13 <= T_2365_13;
    end else begin
      if (T_9487) begin
        if (6'hd == maxDevs_0) begin
          pending_13 <= GEN_0;
        end else begin
          if (gateways_12_valid) begin
            pending_13 <= 1'h1;
          end
        end
      end else begin
        if (gateways_12_valid) begin
          pending_13 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_14 <= T_2365_14;
    end else begin
      if (T_9487) begin
        if (6'he == maxDevs_0) begin
          pending_14 <= GEN_0;
        end else begin
          if (gateways_13_valid) begin
            pending_14 <= 1'h1;
          end
        end
      end else begin
        if (gateways_13_valid) begin
          pending_14 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_15 <= T_2365_15;
    end else begin
      if (T_9487) begin
        if (6'hf == maxDevs_0) begin
          pending_15 <= GEN_0;
        end else begin
          if (gateways_14_valid) begin
            pending_15 <= 1'h1;
          end
        end
      end else begin
        if (gateways_14_valid) begin
          pending_15 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_16 <= T_2365_16;
    end else begin
      if (T_9487) begin
        if (6'h10 == maxDevs_0) begin
          pending_16 <= GEN_0;
        end else begin
          if (gateways_15_valid) begin
            pending_16 <= 1'h1;
          end
        end
      end else begin
        if (gateways_15_valid) begin
          pending_16 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_17 <= T_2365_17;
    end else begin
      if (T_9487) begin
        if (6'h11 == maxDevs_0) begin
          pending_17 <= GEN_0;
        end else begin
          if (gateways_16_valid) begin
            pending_17 <= 1'h1;
          end
        end
      end else begin
        if (gateways_16_valid) begin
          pending_17 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_18 <= T_2365_18;
    end else begin
      if (T_9487) begin
        if (6'h12 == maxDevs_0) begin
          pending_18 <= GEN_0;
        end else begin
          if (gateways_17_valid) begin
            pending_18 <= 1'h1;
          end
        end
      end else begin
        if (gateways_17_valid) begin
          pending_18 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_19 <= T_2365_19;
    end else begin
      if (T_9487) begin
        if (6'h13 == maxDevs_0) begin
          pending_19 <= GEN_0;
        end else begin
          if (gateways_18_valid) begin
            pending_19 <= 1'h1;
          end
        end
      end else begin
        if (gateways_18_valid) begin
          pending_19 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_20 <= T_2365_20;
    end else begin
      if (T_9487) begin
        if (6'h14 == maxDevs_0) begin
          pending_20 <= GEN_0;
        end else begin
          if (gateways_19_valid) begin
            pending_20 <= 1'h1;
          end
        end
      end else begin
        if (gateways_19_valid) begin
          pending_20 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_21 <= T_2365_21;
    end else begin
      if (T_9487) begin
        if (6'h15 == maxDevs_0) begin
          pending_21 <= GEN_0;
        end else begin
          if (gateways_20_valid) begin
            pending_21 <= 1'h1;
          end
        end
      end else begin
        if (gateways_20_valid) begin
          pending_21 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_22 <= T_2365_22;
    end else begin
      if (T_9487) begin
        if (6'h16 == maxDevs_0) begin
          pending_22 <= GEN_0;
        end else begin
          if (gateways_21_valid) begin
            pending_22 <= 1'h1;
          end
        end
      end else begin
        if (gateways_21_valid) begin
          pending_22 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_23 <= T_2365_23;
    end else begin
      if (T_9487) begin
        if (6'h17 == maxDevs_0) begin
          pending_23 <= GEN_0;
        end else begin
          if (gateways_22_valid) begin
            pending_23 <= 1'h1;
          end
        end
      end else begin
        if (gateways_22_valid) begin
          pending_23 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_24 <= T_2365_24;
    end else begin
      if (T_9487) begin
        if (6'h18 == maxDevs_0) begin
          pending_24 <= GEN_0;
        end else begin
          if (gateways_23_valid) begin
            pending_24 <= 1'h1;
          end
        end
      end else begin
        if (gateways_23_valid) begin
          pending_24 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_25 <= T_2365_25;
    end else begin
      if (T_9487) begin
        if (6'h19 == maxDevs_0) begin
          pending_25 <= GEN_0;
        end else begin
          if (gateways_24_valid) begin
            pending_25 <= 1'h1;
          end
        end
      end else begin
        if (gateways_24_valid) begin
          pending_25 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_26 <= T_2365_26;
    end else begin
      if (T_9487) begin
        if (6'h1a == maxDevs_0) begin
          pending_26 <= GEN_0;
        end else begin
          if (gateways_25_valid) begin
            pending_26 <= 1'h1;
          end
        end
      end else begin
        if (gateways_25_valid) begin
          pending_26 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_27 <= T_2365_27;
    end else begin
      if (T_9487) begin
        if (6'h1b == maxDevs_0) begin
          pending_27 <= GEN_0;
        end else begin
          if (gateways_26_valid) begin
            pending_27 <= 1'h1;
          end
        end
      end else begin
        if (gateways_26_valid) begin
          pending_27 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_28 <= T_2365_28;
    end else begin
      if (T_9487) begin
        if (6'h1c == maxDevs_0) begin
          pending_28 <= GEN_0;
        end else begin
          if (gateways_27_valid) begin
            pending_28 <= 1'h1;
          end
        end
      end else begin
        if (gateways_27_valid) begin
          pending_28 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_29 <= T_2365_29;
    end else begin
      if (T_9487) begin
        if (6'h1d == maxDevs_0) begin
          pending_29 <= GEN_0;
        end else begin
          if (gateways_28_valid) begin
            pending_29 <= 1'h1;
          end
        end
      end else begin
        if (gateways_28_valid) begin
          pending_29 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_30 <= T_2365_30;
    end else begin
      if (T_9487) begin
        if (6'h1e == maxDevs_0) begin
          pending_30 <= GEN_0;
        end else begin
          if (gateways_29_valid) begin
            pending_30 <= 1'h1;
          end
        end
      end else begin
        if (gateways_29_valid) begin
          pending_30 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_31 <= T_2365_31;
    end else begin
      if (T_9487) begin
        if (6'h1f == maxDevs_0) begin
          pending_31 <= GEN_0;
        end else begin
          if (gateways_30_valid) begin
            pending_31 <= 1'h1;
          end
        end
      end else begin
        if (gateways_30_valid) begin
          pending_31 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_32 <= T_2365_32;
    end else begin
      if (T_9487) begin
        if (6'h20 == maxDevs_0) begin
          pending_32 <= GEN_0;
        end else begin
          if (gateways_31_valid) begin
            pending_32 <= 1'h1;
          end
        end
      end else begin
        if (gateways_31_valid) begin
          pending_32 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_33 <= T_2365_33;
    end else begin
      if (T_9487) begin
        if (6'h21 == maxDevs_0) begin
          pending_33 <= GEN_0;
        end else begin
          if (gateways_32_valid) begin
            pending_33 <= 1'h1;
          end
        end
      end else begin
        if (gateways_32_valid) begin
          pending_33 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_34 <= T_2365_34;
    end else begin
      if (T_9487) begin
        if (6'h22 == maxDevs_0) begin
          pending_34 <= GEN_0;
        end else begin
          if (gateways_33_valid) begin
            pending_34 <= 1'h1;
          end
        end
      end else begin
        if (gateways_33_valid) begin
          pending_34 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_35 <= T_2365_35;
    end else begin
      if (T_9487) begin
        if (6'h23 == maxDevs_0) begin
          pending_35 <= GEN_0;
        end else begin
          if (gateways_34_valid) begin
            pending_35 <= 1'h1;
          end
        end
      end else begin
        if (gateways_34_valid) begin
          pending_35 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_36 <= T_2365_36;
    end else begin
      if (T_9487) begin
        if (6'h24 == maxDevs_0) begin
          pending_36 <= GEN_0;
        end else begin
          if (gateways_35_valid) begin
            pending_36 <= 1'h1;
          end
        end
      end else begin
        if (gateways_35_valid) begin
          pending_36 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_37 <= T_2365_37;
    end else begin
      if (T_9487) begin
        if (6'h25 == maxDevs_0) begin
          pending_37 <= GEN_0;
        end else begin
          if (gateways_36_valid) begin
            pending_37 <= 1'h1;
          end
        end
      end else begin
        if (gateways_36_valid) begin
          pending_37 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_38 <= T_2365_38;
    end else begin
      if (T_9487) begin
        if (6'h26 == maxDevs_0) begin
          pending_38 <= GEN_0;
        end else begin
          if (gateways_37_valid) begin
            pending_38 <= 1'h1;
          end
        end
      end else begin
        if (gateways_37_valid) begin
          pending_38 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_39 <= T_2365_39;
    end else begin
      if (T_9487) begin
        if (6'h27 == maxDevs_0) begin
          pending_39 <= GEN_0;
        end else begin
          if (gateways_38_valid) begin
            pending_39 <= 1'h1;
          end
        end
      end else begin
        if (gateways_38_valid) begin
          pending_39 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_40 <= T_2365_40;
    end else begin
      if (T_9487) begin
        if (6'h28 == maxDevs_0) begin
          pending_40 <= GEN_0;
        end else begin
          if (gateways_39_valid) begin
            pending_40 <= 1'h1;
          end
        end
      end else begin
        if (gateways_39_valid) begin
          pending_40 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_41 <= T_2365_41;
    end else begin
      if (T_9487) begin
        if (6'h29 == maxDevs_0) begin
          pending_41 <= GEN_0;
        end else begin
          if (gateways_40_valid) begin
            pending_41 <= 1'h1;
          end
        end
      end else begin
        if (gateways_40_valid) begin
          pending_41 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_42 <= T_2365_42;
    end else begin
      if (T_9487) begin
        if (6'h2a == maxDevs_0) begin
          pending_42 <= GEN_0;
        end else begin
          if (gateways_41_valid) begin
            pending_42 <= 1'h1;
          end
        end
      end else begin
        if (gateways_41_valid) begin
          pending_42 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_43 <= T_2365_43;
    end else begin
      if (T_9487) begin
        if (6'h2b == maxDevs_0) begin
          pending_43 <= GEN_0;
        end else begin
          if (gateways_42_valid) begin
            pending_43 <= 1'h1;
          end
        end
      end else begin
        if (gateways_42_valid) begin
          pending_43 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_44 <= T_2365_44;
    end else begin
      if (T_9487) begin
        if (6'h2c == maxDevs_0) begin
          pending_44 <= GEN_0;
        end else begin
          if (gateways_43_valid) begin
            pending_44 <= 1'h1;
          end
        end
      end else begin
        if (gateways_43_valid) begin
          pending_44 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_45 <= T_2365_45;
    end else begin
      if (T_9487) begin
        if (6'h2d == maxDevs_0) begin
          pending_45 <= GEN_0;
        end else begin
          if (gateways_44_valid) begin
            pending_45 <= 1'h1;
          end
        end
      end else begin
        if (gateways_44_valid) begin
          pending_45 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_46 <= T_2365_46;
    end else begin
      if (T_9487) begin
        if (6'h2e == maxDevs_0) begin
          pending_46 <= GEN_0;
        end else begin
          if (gateways_45_valid) begin
            pending_46 <= 1'h1;
          end
        end
      end else begin
        if (gateways_45_valid) begin
          pending_46 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_47 <= T_2365_47;
    end else begin
      if (T_9487) begin
        if (6'h2f == maxDevs_0) begin
          pending_47 <= GEN_0;
        end else begin
          if (gateways_46_valid) begin
            pending_47 <= 1'h1;
          end
        end
      end else begin
        if (gateways_46_valid) begin
          pending_47 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_48 <= T_2365_48;
    end else begin
      if (T_9487) begin
        if (6'h30 == maxDevs_0) begin
          pending_48 <= GEN_0;
        end else begin
          if (gateways_47_valid) begin
            pending_48 <= 1'h1;
          end
        end
      end else begin
        if (gateways_47_valid) begin
          pending_48 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_49 <= T_2365_49;
    end else begin
      if (T_9487) begin
        if (6'h31 == maxDevs_0) begin
          pending_49 <= GEN_0;
        end else begin
          if (gateways_48_valid) begin
            pending_49 <= 1'h1;
          end
        end
      end else begin
        if (gateways_48_valid) begin
          pending_49 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_50 <= T_2365_50;
    end else begin
      if (T_9487) begin
        if (6'h32 == maxDevs_0) begin
          pending_50 <= GEN_0;
        end else begin
          if (gateways_49_valid) begin
            pending_50 <= 1'h1;
          end
        end
      end else begin
        if (gateways_49_valid) begin
          pending_50 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
    if (reset) begin
      pending_51 <= T_2365_51;
    end else begin
      if (T_9487) begin
        if (6'h33 == maxDevs_0) begin
          pending_51 <= GEN_0;
        end else begin
          if (gateways_50_valid) begin
            pending_51 <= 1'h1;
          end
        end
      end else begin
        if (gateways_50_valid) begin
          pending_51 <= 1'h1;
        end
      end
    end
  end

  always @(posedge clock or posedge reset) begin
  if (reset) begin
      enables_0_0 <= 1'h0;
      enables_0_1 <= 1'h0;
      enables_0_2 <= 1'h0;
      enables_0_3 <= 1'h0;
      enables_0_4 <= 1'h0;
      enables_0_5 <= 1'h0;
      enables_0_6 <= 1'h0;
      enables_0_7 <= 1'h0;
      enables_0_8 <= 1'h0;
      enables_0_9 <= 1'h0;
      enables_0_10 <= 1'h0;
      enables_0_11 <= 1'h0;
      enables_0_12 <= 1'h0;
      enables_0_13 <= 1'h0;
      enables_0_14 <= 1'h0;
      enables_0_15 <= 1'h0;
      enables_0_16 <= 1'h0;
      enables_0_17 <= 1'h0;
      enables_0_18 <= 1'h0;
      enables_0_19 <= 1'h0;
      enables_0_20 <= 1'h0;
      enables_0_21 <= 1'h0;
      enables_0_22 <= 1'h0;
      enables_0_23 <= 1'h0;
      enables_0_24 <= 1'h0;
      enables_0_25 <= 1'h0;
      enables_0_26 <= 1'h0;
      enables_0_27 <= 1'h0;
      enables_0_28 <= 1'h0;
      enables_0_29 <= 1'h0;
      enables_0_30 <= 1'h0;
      enables_0_31 <= 1'h0;
      enables_0_32 <= 1'h0;
      enables_0_33 <= 1'h0;
      enables_0_34 <= 1'h0;
      enables_0_35 <= 1'h0;
      enables_0_36 <= 1'h0;
      enables_0_37 <= 1'h0;
      enables_0_38 <= 1'h0;
      enables_0_39 <= 1'h0;
      enables_0_40 <= 1'h0;
      enables_0_41 <= 1'h0;
      enables_0_42 <= 1'h0;
      enables_0_43 <= 1'h0;
      enables_0_44 <= 1'h0;
      enables_0_45 <= 1'h0;
      enables_0_46 <= 1'h0;
      enables_0_47 <= 1'h0;
      enables_0_48 <= 1'h0;
      enables_0_49 <= 1'h0;
      enables_0_50 <= 1'h0;
      enables_0_51 <= 1'h0;
  end
  else begin
    enables_0_0 <= 1'h0;
    if (T_10194) begin
      enables_0_1 <= T_7012;
    end
    if (T_10234) begin
      enables_0_2 <= T_7052;
    end
    if (T_10274) begin
      enables_0_3 <= T_7092;
    end
    if (T_10314) begin
      enables_0_4 <= T_7132;
    end
    if (T_10354) begin
      enables_0_5 <= T_7172;
    end
    if (T_10394) begin
      enables_0_6 <= T_7212;
    end
    if (T_10434) begin
      enables_0_7 <= T_7252;
    end
    if (T_10474) begin
      enables_0_8 <= T_7292;
    end
    if (T_10514) begin
      enables_0_9 <= T_7332;
    end
    if (T_10554) begin
      enables_0_10 <= T_7372;
    end
    if (T_10594) begin
      enables_0_11 <= T_7412;
    end
    if (T_10634) begin
      enables_0_12 <= T_7452;
    end
    if (T_10674) begin
      enables_0_13 <= T_7492;
    end
    if (T_10714) begin
      enables_0_14 <= T_7532;
    end
    if (T_10754) begin
      enables_0_15 <= T_7572;
    end
    if (T_10794) begin
      enables_0_16 <= T_7612;
    end
    if (T_10834) begin
      enables_0_17 <= T_7652;
    end
    if (T_10874) begin
      enables_0_18 <= T_7692;
    end
    if (T_10914) begin
      enables_0_19 <= T_7732;
    end
    if (T_10954) begin
      enables_0_20 <= T_7772;
    end
    if (T_10994) begin
      enables_0_21 <= T_7812;
    end
    if (T_11034) begin
      enables_0_22 <= T_7852;
    end
    if (T_11074) begin
      enables_0_23 <= T_7892;
    end
    if (T_11114) begin
      enables_0_24 <= T_7932;
    end
    if (T_11154) begin
      enables_0_25 <= T_7972;
    end
    if (T_11194) begin
      enables_0_26 <= T_8012;
    end
    if (T_11234) begin
      enables_0_27 <= T_8052;
    end
    if (T_11274) begin
      enables_0_28 <= T_8092;
    end
    if (T_11314) begin
      enables_0_29 <= T_8132;
    end
    if (T_11354) begin
      enables_0_30 <= T_8172;
    end
    if (T_11394) begin
      enables_0_31 <= T_8212;
    end
    if (T_8611) begin
      enables_0_32 <= T_6972;
    end
    if (T_8651) begin
      enables_0_33 <= T_7012;
    end
    if (T_8691) begin
      enables_0_34 <= T_7052;
    end
    if (T_8731) begin
      enables_0_35 <= T_7092;
    end
    if (T_8771) begin
      enables_0_36 <= T_7132;
    end
    if (T_8811) begin
      enables_0_37 <= T_7172;
    end
    if (T_8851) begin
      enables_0_38 <= T_7212;
    end
    if (T_8891) begin
      enables_0_39 <= T_7252;
    end
    if (T_8931) begin
      enables_0_40 <= T_7292;
    end
    if (T_8971) begin
      enables_0_41 <= T_7332;
    end
    if (T_9011) begin
      enables_0_42 <= T_7372;
    end
    if (T_9051) begin
      enables_0_43 <= T_7412;
    end
    if (T_9091) begin
      enables_0_44 <= T_7452;
    end
    if (T_9131) begin
      enables_0_45 <= T_7492;
    end
    if (T_9171) begin
      enables_0_46 <= T_7532;
    end
    if (T_9211) begin
      enables_0_47 <= T_7572;
    end
    if (T_9251) begin
      enables_0_48 <= T_7612;
    end
    if (T_9291) begin
      enables_0_49 <= T_7652;
    end
    if (T_9331) begin
      enables_0_50 <= T_7692;
    end
    if (T_9371) begin
      enables_0_51 <= T_7732;
    end
  end
  end

  always @(posedge clock or posedge reset) begin
  if (reset) begin
      maxDevs_0 <= 6'h0;
  end
  else begin
    if (T_9487) begin
      maxDevs_0 <= 6'h0;
    end else begin
      if (T_3098) begin
        maxDevs_0 <= {{1'd0}, T_2982};
      end else begin
        maxDevs_0 <= T_3101;
      end
    end
  end
  end

  always @(posedge clock or posedge reset) begin
  if (reset) begin
     T_3103 <= 4'h0;
  end
  else begin
    if (T_3098) begin
      if (T_2978) begin
        if (T_2882) begin
          if (T_2834) begin
            if (T_2810) begin
              if (T_2798) begin
                T_3103 <= 4'h8;
              end else begin
                T_3103 <= T_2693;
              end
            end else begin
              if (T_2805) begin
                T_3103 <= T_2695;
              end else begin
                T_3103 <= T_2697;
              end
            end
          end else begin
            if (T_2829) begin
              if (T_2817) begin
                T_3103 <= T_2699;
              end else begin
                T_3103 <= T_2701;
              end
            end else begin
              if (T_2824) begin
                T_3103 <= T_2703;
              end else begin
                T_3103 <= T_2705;
              end
            end
          end
        end else begin
          if (T_2877) begin
            if (T_2853) begin
              if (T_2841) begin
                T_3103 <= T_2707;
              end else begin
                T_3103 <= T_2709;
              end
            end else begin
              if (T_2848) begin
                T_3103 <= T_2711;
              end else begin
                T_3103 <= T_2713;
              end
            end
          end else begin
            if (T_2872) begin
              if (T_2860) begin
                T_3103 <= T_2715;
              end else begin
                T_3103 <= T_2717;
              end
            end else begin
              if (T_2867) begin
                T_3103 <= T_2719;
              end else begin
                T_3103 <= T_2721;
              end
            end
          end
        end
      end else begin
        if (T_2973) begin
          if (T_2925) begin
            if (T_2901) begin
              if (T_2889) begin
                T_3103 <= T_2723;
              end else begin
                T_3103 <= T_2725;
              end
            end else begin
              if (T_2896) begin
                T_3103 <= T_2727;
              end else begin
                T_3103 <= T_2729;
              end
            end
          end else begin
            if (T_2920) begin
              if (T_2908) begin
                T_3103 <= T_2731;
              end else begin
                T_3103 <= T_2733;
              end
            end else begin
              if (T_2915) begin
                T_3103 <= T_2735;
              end else begin
                T_3103 <= T_2737;
              end
            end
          end
        end else begin
          if (T_2968) begin
            if (T_2944) begin
              if (T_2932) begin
                T_3103 <= T_2739;
              end else begin
                T_3103 <= T_2741;
              end
            end else begin
              if (T_2939) begin
                T_3103 <= T_2743;
              end else begin
                T_3103 <= T_2745;
              end
            end
          end else begin
            if (T_2963) begin
              if (T_2951) begin
                T_3103 <= T_2747;
              end else begin
                T_3103 <= T_2749;
              end
            end else begin
              if (T_2958) begin
                T_3103 <= T_2751;
              end else begin
                T_3103 <= T_2753;
              end
            end
          end
        end
      end
    end else begin
      if (T_3093) begin
        if (T_3069) begin
          if (T_3021) begin
            if (T_2997) begin
              if (T_2985) begin
                T_3103 <= T_2755;
              end else begin
                T_3103 <= T_2757;
              end
            end else begin
              if (T_2992) begin
                T_3103 <= T_2759;
              end else begin
                T_3103 <= T_2761;
              end
            end
          end else begin
            if (T_3016) begin
              if (T_3004) begin
                T_3103 <= T_2763;
              end else begin
                T_3103 <= T_2765;
              end
            end else begin
              if (T_3011) begin
                T_3103 <= T_2767;
              end else begin
                T_3103 <= T_2769;
              end
            end
          end
        end else begin
          if (T_3064) begin
            if (T_3040) begin
              if (T_3028) begin
                T_3103 <= T_2771;
              end else begin
                T_3103 <= T_2773;
              end
            end else begin
              if (T_3035) begin
                T_3103 <= T_2775;
              end else begin
                T_3103 <= T_2777;
              end
            end
          end else begin
            if (T_3059) begin
              if (T_3047) begin
                T_3103 <= T_2779;
              end else begin
                T_3103 <= T_2781;
              end
            end else begin
              if (T_3054) begin
                T_3103 <= T_2783;
              end else begin
                T_3103 <= T_2785;
              end
            end
          end
        end
      end else begin
        if (T_3088) begin
          if (T_3076) begin
            T_3103 <= T_2787;
          end else begin
            T_3103 <= T_2789;
          end
        end else begin
          if (T_3083) begin
            T_3103 <= T_2791;
          end else begin
            T_3103 <= T_2793;
          end
        end
      end
    end
  end
  end
endmodule
